* SPICE3 file created from BUFFER_TEST_0.ext - technology: sky130A

.subckt BUFFER_TEST_0 VIN VOUT VSS VDD
X0 VOUT STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X1 VOUT STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VSS STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 VSS STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X4 VOUT STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VOUT STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 VSS STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X7 VOUT STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VSS VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X8 VSS STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 VSS STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VIN VSS VSS sky130_fd_pr__nfet_01v8 ad=0.588 pd=7 as=1.386 ps=16.68 w=0.42 l=0.15
X11 STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VIN VSS VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X12 VSS VIN STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X13 VSS VIN STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X14 STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VIN VSS VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X15 STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VIN VSS VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X16 VSS VIN STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X17 STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VIN VSS VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X18 VSS VIN STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X19 VSS VIN STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VSS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X20 VDD STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.12 as=0.1176 ps=1.12 w=0.84 l=0.15
X21 VOUT STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.12 as=0.1176 ps=1.12 w=0.84 l=0.15
X22 VOUT STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.12 as=0.1176 ps=1.12 w=0.84 l=0.15
X23 VDD STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.2226 pd=2.21 as=0.1176 ps=1.12 w=0.84 l=0.15
X24 VOUT STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.12 as=0.2226 ps=2.21 w=0.84 l=0.15
X25 VDD STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.12 as=0.1176 ps=1.12 w=0.84 l=0.15
X26 VDD STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.12 as=0.1176 ps=1.12 w=0.84 l=0.15
X27 VOUT STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.12 as=0.1176 ps=1.12 w=0.84 l=0.15
X28 VOUT STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.12 as=0.1176 ps=1.12 w=0.84 l=0.15
X29 VDD STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.12 as=0.1176 ps=1.12 w=0.84 l=0.15
X30 VDD VIN STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VDD sky130_fd_pr__pfet_01v8 ad=2.772 pd=26.76 as=1.176 ps=11.2 w=0.84 l=0.15
X31 STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VIN VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X32 STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VIN VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X33 VDD VIN STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X34 STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VIN VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X35 VDD VIN STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X36 VDD VIN STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X37 STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VIN VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X38 STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VIN VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X39 VDD VIN STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
C0 VIN VDD 4.57fF
C1 VOUT VDD 4.42fF
C2 STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VDD 8.38fF
C3 VIN VSS 3.31fF
C4 VDD VSS 14.52fF
C5 VOUT VSS 3.03fF
C6 STAGE2_INV_86799252_PG0_0_0_1677905997_0/li_1179_1411# VSS 7.08fF 
.ends

*=======Added manually========
X1 in out GND VDD BUFFER_TEST_0
V1 VDD GND 1.8
.save i(net1)
V2 in GND pulse(0 1.8 1n 1n 1n 4n 10n)
.save i(in)
**** begin user architecture code

.lib /home/pramit/EDA_TOOLS/skywater-pdk/libraries/sky130_fd_pr/latest/models/sky130.lib.spice tt

.control
save all
tran 1n 20n
plot v(in) v(out)
.endc
