magic
tech sky130A
magscale 1 2
timestamp 1678560175
<< metal1 >>
rect 226 2462 290 2464
rect 226 2410 232 2462
rect 284 2410 290 2462
rect 226 2408 290 2410
rect 312 1622 376 1624
rect 312 1570 318 1622
rect 370 1570 376 1622
rect 312 1568 376 1570
rect 312 1454 376 1456
rect 312 1402 318 1454
rect 370 1402 376 1454
rect 312 1400 376 1402
rect 226 614 290 616
rect 226 562 232 614
rect 284 562 290 614
rect 226 560 290 562
<< via1 >>
rect 232 2410 284 2462
rect 318 1570 370 1622
rect 318 1402 370 1454
rect 232 562 284 614
<< metal2 >>
rect 230 2462 286 2468
rect 230 2410 232 2462
rect 284 2410 286 2462
rect 230 614 286 2410
rect 316 1622 372 1628
rect 316 1570 318 1622
rect 370 1570 372 1622
rect 316 1454 372 1570
rect 316 1402 318 1454
rect 370 1402 372 1454
rect 316 1396 372 1402
rect 230 562 232 614
rect 284 562 286 614
rect 230 556 286 562
use NMOS_S_97312901_X2_Y1_1678559784_1678559786  NMOS_S_97312901_X2_Y1_1678559784_1678559786_0
timestamp 1678560175
transform 1 0 0 0 -1 1512
box 121 56 567 1482
use PMOS_S_78930897_X2_Y1_1678559785_1678559786  PMOS_S_78930897_X2_Y1_1678559785_1678559786_0
timestamp 1678560175
transform 1 0 0 0 1 1512
box 0 0 688 1512
<< end >>
