magic
tech sky130A
magscale 1 2
timestamp 1678552702
<< locali >>
rect 491 1747 499 1781
rect 533 1747 541 1781
rect 1265 1747 1273 1781
rect 1307 1747 1315 1781
rect 491 1613 541 1747
rect 491 1579 499 1613
rect 533 1579 541 1613
rect 663 1579 671 1613
rect 705 1579 713 1613
rect 663 1529 713 1579
rect 663 1495 671 1529
rect 705 1495 713 1529
rect 663 655 671 689
rect 705 655 713 689
rect 663 605 713 655
rect 663 571 671 605
rect 705 571 713 605
<< viali >>
rect 499 1747 533 1781
rect 1273 1747 1307 1781
rect 499 1579 533 1613
rect 671 1579 705 1613
rect 671 1495 705 1529
rect 671 655 705 689
rect 671 571 705 605
<< metal1 >>
rect 312 2882 376 2884
rect 312 2830 318 2882
rect 370 2830 376 2882
rect 312 2828 376 2830
rect 656 2882 720 2884
rect 656 2830 662 2882
rect 714 2830 720 2882
rect 656 2828 720 2830
rect 494 2408 592 2464
rect 482 1781 1324 1792
rect 482 1747 499 1781
rect 533 1747 1273 1781
rect 1307 1747 1324 1781
rect 482 1736 1324 1747
rect 1516 1790 1666 1792
rect 1516 1738 1522 1790
rect 1574 1738 1608 1790
rect 1660 1738 1666 1790
rect 1516 1736 1666 1738
rect 430 1706 806 1708
rect 430 1654 748 1706
rect 800 1654 806 1706
rect 430 1652 806 1654
rect 312 1622 376 1624
rect 312 1570 318 1622
rect 370 1570 376 1622
rect 312 1568 376 1570
rect 482 1613 550 1624
rect 482 1579 499 1613
rect 533 1579 550 1613
rect 482 1568 550 1579
rect 654 1613 722 1624
rect 654 1579 671 1613
rect 705 1579 722 1613
rect 654 1568 722 1579
rect 398 1538 722 1540
rect 398 1486 404 1538
rect 456 1529 722 1538
rect 456 1495 671 1529
rect 705 1495 722 1529
rect 456 1486 722 1495
rect 398 1484 722 1486
rect 742 1454 806 1456
rect 742 1402 748 1454
rect 800 1402 806 1454
rect 742 1400 806 1402
rect 1182 1400 1312 1456
rect 312 1370 376 1372
rect 312 1318 318 1370
rect 370 1318 376 1370
rect 312 1316 376 1318
rect 1430 1286 1580 1288
rect 1430 1234 1436 1286
rect 1488 1234 1522 1286
rect 1574 1234 1580 1286
rect 1430 1232 1580 1234
rect 398 698 722 700
rect 398 646 404 698
rect 456 689 722 698
rect 456 655 671 689
rect 705 655 722 689
rect 456 646 722 655
rect 398 644 722 646
rect 654 605 774 616
rect 654 571 671 605
rect 705 571 774 605
rect 654 560 774 571
rect 140 110 290 112
rect 140 58 146 110
rect 198 58 232 110
rect 284 58 290 110
rect 140 56 290 58
<< via1 >>
rect 318 2830 370 2882
rect 662 2830 714 2882
rect 1522 1738 1574 1790
rect 1608 1738 1660 1790
rect 748 1654 800 1706
rect 318 1570 370 1622
rect 404 1486 456 1538
rect 748 1402 800 1454
rect 318 1318 370 1370
rect 1436 1234 1488 1286
rect 1522 1234 1574 1286
rect 404 646 456 698
rect 146 58 198 110
rect 232 58 284 110
<< metal2 >>
rect 316 2882 372 2888
rect 316 2830 318 2882
rect 370 2830 372 2882
rect 316 1792 372 2830
rect 316 1727 372 1736
rect 660 2882 716 2888
rect 660 2830 662 2882
rect 714 2830 716 2882
rect 660 1792 716 2830
rect 660 1727 716 1736
rect 1004 1792 1060 1801
rect 746 1706 802 1712
rect 746 1654 748 1706
rect 800 1654 802 1706
rect 316 1622 372 1628
rect 316 1570 318 1622
rect 370 1570 372 1622
rect 316 1370 372 1570
rect 402 1538 458 1544
rect 402 1486 404 1538
rect 456 1486 458 1538
rect 402 1428 458 1486
rect 746 1454 802 1654
rect 746 1402 748 1454
rect 800 1402 802 1454
rect 746 1396 802 1402
rect 316 1318 318 1370
rect 370 1318 372 1370
rect 1004 1344 1060 1736
rect 1434 1792 1490 1801
rect 316 1312 372 1318
rect 1434 1286 1490 1736
rect 1520 1790 1576 1796
rect 1520 1738 1522 1790
rect 1574 1738 1576 1790
rect 1520 1732 1576 1738
rect 1606 1790 1662 1796
rect 1606 1738 1608 1790
rect 1660 1738 1662 1790
rect 1434 1234 1436 1286
rect 1488 1234 1490 1286
rect 1434 1228 1490 1234
rect 1520 1286 1576 1292
rect 1520 1234 1522 1286
rect 1574 1234 1576 1286
rect 1520 1228 1576 1234
rect 402 698 458 704
rect 402 646 404 698
rect 456 646 458 698
rect 402 640 458 646
rect 144 110 200 116
rect 144 58 146 110
rect 198 58 200 110
rect 144 28 200 58
rect 230 110 286 168
rect 230 58 232 110
rect 284 58 286 110
rect 230 52 286 58
rect 144 -37 200 -28
rect 1606 28 1662 1738
rect 1606 -37 1662 -28
<< via2 >>
rect 316 1736 372 1792
rect 660 1736 716 1792
rect 1004 1736 1060 1792
rect 1434 1736 1490 1792
rect 144 -28 200 28
rect 1606 -28 1662 28
<< metal3 >>
rect -80 1796 2448 1844
rect -80 1792 2336 1796
rect -80 1736 316 1792
rect 372 1736 660 1792
rect 716 1736 1004 1792
rect 1060 1736 1434 1792
rect 1490 1736 2336 1792
rect -80 1732 2336 1736
rect 2400 1732 2448 1796
rect -80 1684 2448 1732
rect -80 32 2448 80
rect -80 -32 -32 32
rect 32 28 2448 32
rect 32 -28 144 28
rect 200 -28 1606 28
rect 1662 -28 2448 28
rect 32 -32 2448 -28
rect -80 -80 2448 -32
<< via3 >>
rect 2336 1732 2400 1796
rect -32 -32 32 32
<< metal4 >>
rect -118 32 118 1882
rect -118 -32 -32 32
rect 32 -32 118 32
rect -118 -118 118 -32
rect 2250 1796 2486 1882
rect 2250 1732 2336 1796
rect 2400 1732 2486 1796
rect 2250 -118 2486 1732
use INV_14817437_PG0_0_0_1678552160  INV_14817437_PG0_0_0_1678552160_0
timestamp 1678552702
transform 1 0 1204 0 1 0
box 0 30 516 3024
use NMOS_4T_90354340_X1_Y1_1678552161  NMOS_4T_90354340_X1_Y1_1678552161_0
timestamp 1678552702
transform 1 0 602 0 1 1512
box 52 56 395 1482
use NMOS_4T_90354340_X1_Y1_1678552161  NMOS_4T_90354340_X1_Y1_1678552161_1
timestamp 1678552702
transform -1 0 602 0 1 1512
box 52 56 395 1482
use NMOS_S_25628869_X1_Y1_1678552162  NMOS_S_25628869_X1_Y1_1678552162_0
timestamp 1678552702
transform 1 0 688 0 -1 1512
box 52 56 395 1482
use SCM_PMOS_73046675_X1_Y1_1678552163  SCM_PMOS_73046675_X1_Y1_1678552163_0
timestamp 1678552702
transform -1 0 688 0 -1 1512
box 0 0 688 1512
<< labels >>
flabel metal1 s 774 2436 774 2436 0 FreeSerif 0 0 0 0 INN
port 1 nsew
flabel metal2 s 1032 1554 1032 1554 0 FreeSerif 0 0 0 0 GND
port 2 nsew
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
port 2 nsew
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
port 2 nsew
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
port 2 nsew
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
port 2 nsew
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
port 2 nsew
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
port 2 nsew
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
port 2 nsew
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
port 2 nsew
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
port 2 nsew
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
port 2 nsew
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
port 2 nsew
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
port 2 nsew
flabel metal2 s 258 126 258 126 0 FreeSerif 0 0 0 0 VDD
port 3 nsew
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VDD
port 3 nsew
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VDD
port 3 nsew
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VDD
port 3 nsew
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VDD
port 3 nsew
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VDD
port 3 nsew
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VDD
port 3 nsew
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VDD
port 3 nsew
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VDD
port 3 nsew
flabel metal1 s 1206 1430 1206 1430 1 FreeSans 480 0 0 0 OUT
port 4 n
flabel metal1 s 566 2430 566 2430 1 FreeSans 480 0 0 0 INP
port 5 n
<< end >>
