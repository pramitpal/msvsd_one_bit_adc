magic
tech sky130A
magscale 1 2
timestamp 1678560175
<< pwell >>
rect 215 1206 473 1482
rect 121 457 567 677
<< nmos >>
rect 200 483 230 651
rect 286 483 316 651
rect 372 483 402 651
rect 458 483 488 651
<< ndiff >>
rect 147 601 200 651
rect 147 567 155 601
rect 189 567 200 601
rect 147 533 200 567
rect 147 499 155 533
rect 189 499 200 533
rect 147 483 200 499
rect 230 601 286 651
rect 230 567 241 601
rect 275 567 286 601
rect 230 533 286 567
rect 230 499 241 533
rect 275 499 286 533
rect 230 483 286 499
rect 316 601 372 651
rect 316 567 327 601
rect 361 567 372 601
rect 316 533 372 567
rect 316 499 327 533
rect 361 499 372 533
rect 316 483 372 499
rect 402 601 458 651
rect 402 567 413 601
rect 447 567 458 601
rect 402 533 458 567
rect 402 499 413 533
rect 447 499 458 533
rect 402 483 458 499
rect 488 601 541 651
rect 488 567 499 601
rect 533 567 541 601
rect 488 533 541 567
rect 488 499 499 533
rect 533 499 541 533
rect 488 483 541 499
<< ndiffc >>
rect 155 567 189 601
rect 155 499 189 533
rect 241 567 275 601
rect 241 499 275 533
rect 327 567 361 601
rect 327 499 361 533
rect 413 567 447 601
rect 413 499 447 533
rect 499 567 533 601
rect 499 499 533 533
<< psubdiff >>
rect 241 1361 275 1456
rect 241 1232 275 1327
rect 413 1361 447 1456
rect 413 1232 447 1327
<< psubdiffcont >>
rect 241 1327 275 1361
rect 413 1327 447 1361
<< poly >>
rect 200 941 316 951
rect 200 907 241 941
rect 275 907 316 941
rect 200 897 316 907
rect 200 651 230 897
rect 286 651 316 897
rect 372 941 488 951
rect 372 907 413 941
rect 447 907 488 941
rect 372 897 488 907
rect 372 651 402 897
rect 458 651 488 897
rect 200 252 230 483
rect 286 252 316 483
rect 372 252 402 483
rect 458 252 488 483
<< polycont >>
rect 241 907 275 941
rect 413 907 447 941
<< locali >>
rect 233 1361 283 1445
rect 233 1327 241 1361
rect 275 1327 283 1361
rect 233 1243 283 1327
rect 405 1361 455 1445
rect 405 1327 413 1361
rect 447 1327 455 1361
rect 405 1243 455 1327
rect 233 941 283 1025
rect 233 907 241 941
rect 275 907 283 941
rect 233 823 283 907
rect 405 941 455 1025
rect 405 907 413 941
rect 447 907 455 941
rect 405 823 455 907
rect 147 601 197 773
rect 147 567 155 601
rect 189 567 197 601
rect 147 533 197 567
rect 147 499 155 533
rect 189 499 197 533
rect 147 185 197 499
rect 147 151 155 185
rect 189 151 197 185
rect 147 67 197 151
rect 233 601 283 773
rect 233 567 241 601
rect 275 567 283 601
rect 233 533 283 567
rect 233 499 241 533
rect 275 499 283 533
rect 233 101 283 499
rect 233 67 241 101
rect 275 67 283 101
rect 319 601 369 773
rect 319 567 327 601
rect 361 567 369 601
rect 319 533 369 567
rect 319 499 327 533
rect 361 499 369 533
rect 319 185 369 499
rect 319 151 327 185
rect 361 151 369 185
rect 319 67 369 151
rect 405 601 455 773
rect 405 567 413 601
rect 447 567 455 601
rect 405 533 455 567
rect 405 499 413 533
rect 447 499 455 533
rect 405 101 455 499
rect 405 67 413 101
rect 447 67 455 101
rect 491 601 541 773
rect 491 567 499 601
rect 533 567 541 601
rect 491 533 541 567
rect 491 499 499 533
rect 533 499 541 533
rect 491 185 541 499
rect 491 151 499 185
rect 533 151 541 185
rect 491 67 541 151
<< viali >>
rect 241 1327 275 1361
rect 413 1327 447 1361
rect 241 907 275 941
rect 413 907 447 941
rect 155 151 189 185
rect 241 67 275 101
rect 327 151 361 185
rect 413 67 447 101
rect 499 151 533 185
<< metal1 >>
rect 224 1361 464 1372
rect 224 1327 241 1361
rect 275 1327 413 1361
rect 447 1327 464 1361
rect 224 1316 464 1327
rect 224 941 464 952
rect 224 907 241 941
rect 275 907 413 941
rect 447 907 464 941
rect 224 896 464 907
rect 138 185 550 196
rect 138 151 155 185
rect 189 151 327 185
rect 361 151 499 185
rect 533 151 550 185
rect 138 140 550 151
rect 224 101 464 112
rect 224 67 241 101
rect 275 67 413 101
rect 447 67 464 101
rect 224 56 464 67
<< end >>
