* SPICE3 file created from adc.ext - technology: sky130A

.subckt adc INP GND VDD INN OUT
X0 GND INP sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X1 GND m3_4894_4713# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X2 GND li_577_5947# OUT GND sky130_fd_pr__nfet_01v8 ad=0.2226 pd=2.21 as=0.1176 ps=1.12 w=0.84 l=0.15
X3 OUT li_577_5947# GND GND sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2226 ps=2.21 w=0.84 l=0.15
X4 GND li_577_5947# OUT GND sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.1176 ps=1.12 w=0.84 l=0.15
X5 OUT li_577_5947# GND GND sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.1176 ps=1.12 w=0.84 l=0.15
X6 OUT li_577_5947# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.12 as=0.2226 ps=2.21 w=0.84 l=0.15
X7 VDD li_577_5947# OUT VDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.12 as=0.1176 ps=1.12 w=0.84 l=0.15
X8 OUT li_577_5947# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.12 as=0.1176 ps=1.12 w=0.84 l=0.15
X9 VDD li_577_5947# OUT VDD sky130_fd_pr__pfet_01v8 ad=0.2226 pd=2.21 as=0.1176 ps=1.12 w=0.84 l=0.15
X10 GND m3_4464_2589# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X11 GND INP m3_4464_2589# GND sky130_fd_pr__nfet_01v8 ad=0.2226 pd=2.21 as=0.1176 ps=1.12 w=0.84 l=0.15
X12 m3_4464_2589# INP GND GND sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2226 ps=2.21 w=0.84 l=0.15
X13 GND INP m3_4464_2589# GND sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.1176 ps=1.12 w=0.84 l=0.15
X14 m3_4464_2589# INP GND GND sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.1176 ps=1.12 w=0.84 l=0.15
X15 m3_4464_2589# INP VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.12 as=0.2226 ps=2.21 w=0.84 l=0.15
X16 VDD INP m3_4464_2589# VDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.12 as=0.1176 ps=1.12 w=0.84 l=0.15
X17 m3_4464_2589# INP VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.12 as=0.1176 ps=1.12 w=0.84 l=0.15
X18 VDD INP m3_4464_2589# VDD sky130_fd_pr__pfet_01v8 ad=0.2226 pd=2.21 as=0.1176 ps=1.12 w=0.84 l=0.15
X19 GND m1_1258_5936# m1_1860_5852# GND sky130_fd_pr__nfet_01v8 ad=0.2226 pd=2.21 as=0.1176 ps=1.12 w=0.84 l=0.15
X20 m1_1860_5852# m1_1258_5936# GND GND sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2226 ps=2.21 w=0.84 l=0.15
X21 GND m1_1258_5936# m1_1860_5852# GND sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.1176 ps=1.12 w=0.84 l=0.15
X22 m1_1860_5852# m1_1258_5936# GND GND sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.1176 ps=1.12 w=0.84 l=0.15
X23 INP m3_4894_4713# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.12 as=0.2226 ps=2.21 w=0.84 l=0.15
X24 VDD m3_4894_4713# INP VDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.12 as=0.1176 ps=1.12 w=0.84 l=0.15
X25 INP m3_4894_4713# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.12 as=0.1176 ps=1.12 w=0.84 l=0.15
X26 VDD m3_4894_4713# INP VDD sky130_fd_pr__pfet_01v8 ad=0.2226 pd=2.21 as=0.1176 ps=1.12 w=0.84 l=0.15
X27 GND m3_4894_4713# INP GND sky130_fd_pr__nfet_01v8 ad=3.402 pd=33.3 as=0.4704 ps=4.48 w=0.84 l=0.15
X28 INP m3_4894_4713# GND GND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X29 GND m3_4894_4713# INP GND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X30 INP m3_4894_4713# GND GND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X31 m3_4894_4713# m3_4464_2589# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.4704 pd=4.48 as=3.8724 ps=37.78 w=0.84 l=0.15
X32 VDD m3_4464_2589# m3_4894_4713# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X33 m3_4894_4713# m3_4464_2589# VDD VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X34 VDD m3_4464_2589# m3_4894_4713# VDD sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X35 GND m3_4464_2589# m3_4894_4713# GND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.4704 ps=4.48 w=0.84 l=0.15
X36 m3_4894_4713# m3_4464_2589# GND GND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X37 GND m3_4464_2589# m3_4894_4713# GND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X38 m3_4894_4713# m3_4464_2589# GND GND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X39 VDD m1_1258_5936# m1_1258_5936# VDD sky130_fd_pr__pfet_01v8 ad=0.2226 pd=2.21 as=0.1176 ps=1.12 w=0.84 l=0.15
X40 li_577_5947# m1_1258_5936# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.12 as=0.1176 ps=1.12 w=0.84 l=0.15
X41 m1_1258_5936# m1_1258_5936# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.12 as=0.2226 ps=2.21 w=0.84 l=0.15
X42 VDD m1_1258_5936# m1_1258_5936# VDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.12 as=0.1176 ps=1.12 w=0.84 l=0.15
X43 VDD m1_1258_5936# li_577_5947# VDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.12 as=0.1176 ps=1.12 w=0.84 l=0.15
X44 li_577_5947# m1_1258_5936# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.12 as=0.1176 ps=1.12 w=0.84 l=0.15
X45 m1_1258_5936# m1_1258_5936# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.12 as=0.1176 ps=1.12 w=0.84 l=0.15
X46 VDD m1_1258_5936# li_577_5947# VDD sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.12 as=0.1176 ps=1.12 w=0.84 l=0.15
X47 m1_1860_5852# INN m1_1258_5936# GND sky130_fd_pr__nfet_01v8 ad=0.2226 pd=2.21 as=0.1176 ps=1.12 w=0.84 l=0.15
X48 m1_1258_5936# INN m1_1860_5852# GND sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2226 ps=2.21 w=0.84 l=0.15
X49 m1_1860_5852# INN m1_1258_5936# GND sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.1176 ps=1.12 w=0.84 l=0.15
X50 m1_1258_5936# INN m1_1860_5852# GND sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.1176 ps=1.12 w=0.84 l=0.15
X51 m1_1860_5852# INP li_577_5947# GND sky130_fd_pr__nfet_01v8 ad=1.8312 pd=17.8 as=0.4704 ps=4.48 w=0.84 l=0.15
X52 li_577_5947# INP m1_1860_5852# GND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X53 m1_1860_5852# INP li_577_5947# GND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X54 li_577_5947# INP m1_1860_5852# GND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
C0 VDD m3_4464_2589# 5.36fF
C1 VDD INP 5.02fF
C2 VDD m1_1258_5936# 5.23fF
C3 m3_4894_4713# VDD 4.40fF
C4 VDD li_577_5947# 3.87fF
C5 m3_4464_2589# GND 7.43fF 
C6 INP GND 10.39fF
C7 m3_4894_4713# GND 6.90fF 
C8 m1_1860_5852# GND 2.04fF 
C9 VDD GND 22.06fF
.ends


x1 INP GND VDD INN OUT adc

V1 VDD GND 1.8
.save i(v1)
V2 INN GND 1
.save i(v2)

.lib /home/pramit/EDA_TOOLS/skywater-pdk/libraries/sky130_fd_pr/latest/models/sky130.lib.spice tt



.tran 0.1n 25n
.save all
.control

run
plot INP INN OUT
.endc
.end
