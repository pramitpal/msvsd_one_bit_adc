magic
tech sky130A
magscale 1 2
timestamp 1678197492
<< viali >>
rect 5181 9129 5215 9163
rect 3985 9061 4019 9095
rect 2053 8993 2087 9027
rect 2329 8925 2363 8959
rect 4169 8925 4203 8959
rect 4261 8925 4295 8959
rect 4997 8925 5031 8959
rect 3985 8857 4019 8891
rect 1685 8585 1719 8619
rect 5181 8585 5215 8619
rect 1869 8449 1903 8483
rect 4997 8449 5031 8483
rect 3525 7293 3559 7327
rect 3801 7293 3835 7327
rect 5273 7157 5307 7191
rect 2329 6817 2363 6851
rect 4905 6817 4939 6851
rect 2697 6749 2731 6783
rect 4997 6749 5031 6783
rect 2605 6681 2639 6715
rect 2513 6613 2547 6647
rect 2881 6613 2915 6647
rect 2053 6273 2087 6307
rect 2605 6273 2639 6307
rect 5181 6273 5215 6307
rect 4997 6137 5031 6171
rect 1961 6069 1995 6103
rect 3893 6069 3927 6103
rect 3433 5797 3467 5831
rect 3157 5729 3191 5763
rect 1869 5661 1903 5695
rect 2053 5661 2087 5695
rect 3065 5661 3099 5695
rect 5181 5661 5215 5695
rect 5089 5593 5123 5627
rect 1961 5525 1995 5559
rect 4261 5321 4295 5355
rect 2221 5253 2255 5287
rect 2421 5253 2455 5287
rect 2973 5185 3007 5219
rect 2053 5049 2087 5083
rect 2237 4981 2271 5015
rect 4077 4777 4111 4811
rect 2421 4709 2455 4743
rect 1869 4573 1903 4607
rect 2605 4573 2639 4607
rect 3157 4573 3191 4607
rect 3985 4573 4019 4607
rect 4813 4573 4847 4607
rect 1685 4437 1719 4471
rect 3341 4437 3375 4471
rect 4721 4437 4755 4471
rect 1777 4097 1811 4131
rect 4629 4097 4663 4131
rect 4721 4097 4755 4131
rect 1685 4029 1719 4063
rect 2237 4029 2271 4063
rect 2513 4029 2547 4063
rect 3985 3893 4019 3927
rect 1685 3689 1719 3723
rect 3433 3485 3467 3519
rect 4169 3485 4203 3519
rect 4813 3485 4847 3519
rect 5089 3485 5123 3519
rect 5273 3485 5307 3519
rect 3157 3417 3191 3451
rect 4629 3417 4663 3451
rect 4077 3349 4111 3383
rect 5273 3145 5307 3179
rect 3801 3077 3835 3111
rect 2237 3009 2271 3043
rect 2329 2941 2363 2975
rect 2605 2941 2639 2975
rect 3525 2941 3559 2975
rect 2145 2601 2179 2635
rect 5181 2601 5215 2635
rect 3433 2397 3467 2431
rect 4537 2397 4571 2431
rect 4997 2397 5031 2431
rect 4353 2261 4387 2295
<< metal1 >>
rect 1104 9274 5796 9296
rect 1104 9222 1950 9274
rect 2002 9222 2014 9274
rect 2066 9222 2078 9274
rect 2130 9222 2142 9274
rect 2194 9222 2206 9274
rect 2258 9222 5796 9274
rect 1104 9200 5796 9222
rect 5166 9120 5172 9172
rect 5224 9120 5230 9172
rect 2958 9052 2964 9104
rect 3016 9092 3022 9104
rect 3973 9095 4031 9101
rect 3973 9092 3985 9095
rect 3016 9064 3985 9092
rect 3016 9052 3022 9064
rect 3973 9061 3985 9064
rect 4019 9061 4031 9095
rect 3973 9055 4031 9061
rect 1854 8984 1860 9036
rect 1912 9024 1918 9036
rect 2041 9027 2099 9033
rect 2041 9024 2053 9027
rect 1912 8996 2053 9024
rect 1912 8984 1918 8996
rect 2041 8993 2053 8996
rect 2087 8993 2099 9027
rect 2041 8987 2099 8993
rect 2317 8959 2375 8965
rect 2317 8925 2329 8959
rect 2363 8956 2375 8959
rect 2406 8956 2412 8968
rect 2363 8928 2412 8956
rect 2363 8925 2375 8928
rect 2317 8919 2375 8925
rect 2406 8916 2412 8928
rect 2464 8956 2470 8968
rect 4157 8959 4215 8965
rect 4157 8956 4169 8959
rect 2464 8928 4169 8956
rect 2464 8916 2470 8928
rect 4157 8925 4169 8928
rect 4203 8925 4215 8959
rect 4157 8919 4215 8925
rect 4246 8916 4252 8968
rect 4304 8916 4310 8968
rect 4338 8916 4344 8968
rect 4396 8956 4402 8968
rect 4985 8959 5043 8965
rect 4985 8956 4997 8959
rect 4396 8928 4997 8956
rect 4396 8916 4402 8928
rect 4985 8925 4997 8928
rect 5031 8925 5043 8959
rect 4985 8919 5043 8925
rect 3050 8848 3056 8900
rect 3108 8888 3114 8900
rect 3973 8891 4031 8897
rect 3973 8888 3985 8891
rect 3108 8860 3985 8888
rect 3108 8848 3114 8860
rect 3973 8857 3985 8860
rect 4019 8857 4031 8891
rect 3973 8851 4031 8857
rect 1104 8730 5796 8752
rect 1104 8678 2610 8730
rect 2662 8678 2674 8730
rect 2726 8678 2738 8730
rect 2790 8678 2802 8730
rect 2854 8678 2866 8730
rect 2918 8678 5796 8730
rect 1104 8656 5796 8678
rect 934 8576 940 8628
rect 992 8616 998 8628
rect 1673 8619 1731 8625
rect 1673 8616 1685 8619
rect 992 8588 1685 8616
rect 992 8576 998 8588
rect 1673 8585 1685 8588
rect 1719 8585 1731 8619
rect 1673 8579 1731 8585
rect 5169 8619 5227 8625
rect 5169 8585 5181 8619
rect 5215 8616 5227 8619
rect 5902 8616 5908 8628
rect 5215 8588 5908 8616
rect 5215 8585 5227 8588
rect 5169 8579 5227 8585
rect 5902 8576 5908 8588
rect 5960 8576 5966 8628
rect 1857 8483 1915 8489
rect 1857 8449 1869 8483
rect 1903 8480 1915 8483
rect 2498 8480 2504 8492
rect 1903 8452 2504 8480
rect 1903 8449 1915 8452
rect 1857 8443 1915 8449
rect 2498 8440 2504 8452
rect 2556 8440 2562 8492
rect 4982 8440 4988 8492
rect 5040 8440 5046 8492
rect 1104 8186 5796 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 5796 8186
rect 1104 8112 5796 8134
rect 1104 7642 5796 7664
rect 1104 7590 2610 7642
rect 2662 7590 2674 7642
rect 2726 7590 2738 7642
rect 2790 7590 2802 7642
rect 2854 7590 2866 7642
rect 2918 7590 5796 7642
rect 1104 7568 5796 7590
rect 4890 7352 4896 7404
rect 4948 7352 4954 7404
rect 3513 7327 3571 7333
rect 3513 7293 3525 7327
rect 3559 7293 3571 7327
rect 3513 7287 3571 7293
rect 3528 7188 3556 7287
rect 3786 7284 3792 7336
rect 3844 7284 3850 7336
rect 3878 7188 3884 7200
rect 3528 7160 3884 7188
rect 3878 7148 3884 7160
rect 3936 7148 3942 7200
rect 5258 7148 5264 7200
rect 5316 7148 5322 7200
rect 1104 7098 5796 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 5796 7098
rect 1104 7024 5796 7046
rect 1762 6808 1768 6860
rect 1820 6848 1826 6860
rect 2317 6851 2375 6857
rect 2317 6848 2329 6851
rect 1820 6820 2329 6848
rect 1820 6808 1826 6820
rect 2317 6817 2329 6820
rect 2363 6848 2375 6851
rect 4338 6848 4344 6860
rect 2363 6820 4344 6848
rect 2363 6817 2375 6820
rect 2317 6811 2375 6817
rect 4338 6808 4344 6820
rect 4396 6808 4402 6860
rect 4890 6808 4896 6860
rect 4948 6808 4954 6860
rect 2222 6740 2228 6792
rect 2280 6780 2286 6792
rect 2685 6783 2743 6789
rect 2685 6780 2697 6783
rect 2280 6752 2697 6780
rect 2280 6740 2286 6752
rect 2685 6749 2697 6752
rect 2731 6780 2743 6783
rect 4246 6780 4252 6792
rect 2731 6752 4252 6780
rect 2731 6749 2743 6752
rect 2685 6743 2743 6749
rect 4246 6740 4252 6752
rect 4304 6740 4310 6792
rect 4706 6740 4712 6792
rect 4764 6780 4770 6792
rect 4985 6783 5043 6789
rect 4985 6780 4997 6783
rect 4764 6752 4997 6780
rect 4764 6740 4770 6752
rect 4985 6749 4997 6752
rect 5031 6749 5043 6783
rect 4985 6743 5043 6749
rect 2593 6715 2651 6721
rect 2593 6681 2605 6715
rect 2639 6712 2651 6715
rect 3050 6712 3056 6724
rect 2639 6684 3056 6712
rect 2639 6681 2651 6684
rect 2593 6675 2651 6681
rect 3050 6672 3056 6684
rect 3108 6672 3114 6724
rect 2406 6604 2412 6656
rect 2464 6644 2470 6656
rect 2501 6647 2559 6653
rect 2501 6644 2513 6647
rect 2464 6616 2513 6644
rect 2464 6604 2470 6616
rect 2501 6613 2513 6616
rect 2547 6613 2559 6647
rect 2501 6607 2559 6613
rect 2869 6647 2927 6653
rect 2869 6613 2881 6647
rect 2915 6644 2927 6647
rect 4154 6644 4160 6656
rect 2915 6616 4160 6644
rect 2915 6613 2927 6616
rect 2869 6607 2927 6613
rect 4154 6604 4160 6616
rect 4212 6604 4218 6656
rect 1104 6554 5796 6576
rect 1104 6502 2610 6554
rect 2662 6502 2674 6554
rect 2726 6502 2738 6554
rect 2790 6502 2802 6554
rect 2854 6502 2866 6554
rect 2918 6502 5796 6554
rect 1104 6480 5796 6502
rect 2041 6307 2099 6313
rect 2041 6273 2053 6307
rect 2087 6304 2099 6307
rect 2314 6304 2320 6316
rect 2087 6276 2320 6304
rect 2087 6273 2099 6276
rect 2041 6267 2099 6273
rect 2314 6264 2320 6276
rect 2372 6264 2378 6316
rect 2593 6307 2651 6313
rect 2593 6273 2605 6307
rect 2639 6304 2651 6307
rect 4062 6304 4068 6316
rect 2639 6276 4068 6304
rect 2639 6273 2651 6276
rect 2593 6267 2651 6273
rect 4062 6264 4068 6276
rect 4120 6264 4126 6316
rect 5169 6307 5227 6313
rect 5169 6273 5181 6307
rect 5215 6304 5227 6307
rect 5902 6304 5908 6316
rect 5215 6276 5908 6304
rect 5215 6273 5227 6276
rect 5169 6267 5227 6273
rect 5902 6264 5908 6276
rect 5960 6264 5966 6316
rect 4706 6128 4712 6180
rect 4764 6168 4770 6180
rect 4985 6171 5043 6177
rect 4985 6168 4997 6171
rect 4764 6140 4997 6168
rect 4764 6128 4770 6140
rect 4985 6137 4997 6140
rect 5031 6137 5043 6171
rect 4985 6131 5043 6137
rect 1854 6060 1860 6112
rect 1912 6100 1918 6112
rect 1949 6103 2007 6109
rect 1949 6100 1961 6103
rect 1912 6072 1961 6100
rect 1912 6060 1918 6072
rect 1949 6069 1961 6072
rect 1995 6069 2007 6103
rect 1949 6063 2007 6069
rect 3878 6060 3884 6112
rect 3936 6060 3942 6112
rect 1104 6010 5796 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 5796 6010
rect 1104 5936 5796 5958
rect 3421 5831 3479 5837
rect 3421 5797 3433 5831
rect 3467 5828 3479 5831
rect 3786 5828 3792 5840
rect 3467 5800 3792 5828
rect 3467 5797 3479 5800
rect 3421 5791 3479 5797
rect 3786 5788 3792 5800
rect 3844 5788 3850 5840
rect 2498 5720 2504 5772
rect 2556 5760 2562 5772
rect 3145 5763 3203 5769
rect 2556 5732 3096 5760
rect 2556 5720 2562 5732
rect 1857 5695 1915 5701
rect 1857 5661 1869 5695
rect 1903 5692 1915 5695
rect 1946 5692 1952 5704
rect 1903 5664 1952 5692
rect 1903 5661 1915 5664
rect 1857 5655 1915 5661
rect 1946 5652 1952 5664
rect 2004 5652 2010 5704
rect 2041 5695 2099 5701
rect 2041 5661 2053 5695
rect 2087 5692 2099 5695
rect 2866 5692 2872 5704
rect 2087 5664 2872 5692
rect 2087 5661 2099 5664
rect 2041 5655 2099 5661
rect 2866 5652 2872 5664
rect 2924 5652 2930 5704
rect 3068 5701 3096 5732
rect 3145 5729 3157 5763
rect 3191 5760 3203 5763
rect 4154 5760 4160 5772
rect 3191 5732 4160 5760
rect 3191 5729 3203 5732
rect 3145 5723 3203 5729
rect 4154 5720 4160 5732
rect 4212 5760 4218 5772
rect 4798 5760 4804 5772
rect 4212 5732 4804 5760
rect 4212 5720 4218 5732
rect 4798 5720 4804 5732
rect 4856 5720 4862 5772
rect 3053 5695 3111 5701
rect 3053 5661 3065 5695
rect 3099 5661 3111 5695
rect 3053 5655 3111 5661
rect 3068 5624 3096 5655
rect 4522 5652 4528 5704
rect 4580 5692 4586 5704
rect 5169 5695 5227 5701
rect 5169 5692 5181 5695
rect 4580 5664 5181 5692
rect 4580 5652 4586 5664
rect 5169 5661 5181 5664
rect 5215 5692 5227 5695
rect 5258 5692 5264 5704
rect 5215 5664 5264 5692
rect 5215 5661 5227 5664
rect 5169 5655 5227 5661
rect 5258 5652 5264 5664
rect 5316 5652 5322 5704
rect 5077 5627 5135 5633
rect 5077 5624 5089 5627
rect 3068 5596 5089 5624
rect 5077 5593 5089 5596
rect 5123 5593 5135 5627
rect 5077 5587 5135 5593
rect 1949 5559 2007 5565
rect 1949 5525 1961 5559
rect 1995 5556 2007 5559
rect 3786 5556 3792 5568
rect 1995 5528 3792 5556
rect 1995 5525 2007 5528
rect 1949 5519 2007 5525
rect 3786 5516 3792 5528
rect 3844 5516 3850 5568
rect 1104 5466 5796 5488
rect 1104 5414 2610 5466
rect 2662 5414 2674 5466
rect 2726 5414 2738 5466
rect 2790 5414 2802 5466
rect 2854 5414 2866 5466
rect 2918 5414 5796 5466
rect 1104 5392 5796 5414
rect 4062 5312 4068 5364
rect 4120 5352 4126 5364
rect 4249 5355 4307 5361
rect 4249 5352 4261 5355
rect 4120 5324 4261 5352
rect 4120 5312 4126 5324
rect 4249 5321 4261 5324
rect 4295 5321 4307 5355
rect 4249 5315 4307 5321
rect 2209 5287 2267 5293
rect 2209 5253 2221 5287
rect 2255 5284 2267 5287
rect 2314 5284 2320 5296
rect 2255 5256 2320 5284
rect 2255 5253 2267 5256
rect 2209 5247 2267 5253
rect 2314 5244 2320 5256
rect 2372 5244 2378 5296
rect 2406 5244 2412 5296
rect 2464 5244 2470 5296
rect 934 5176 940 5228
rect 992 5216 998 5228
rect 2961 5219 3019 5225
rect 2961 5216 2973 5219
rect 992 5188 2973 5216
rect 992 5176 998 5188
rect 2961 5185 2973 5188
rect 3007 5185 3019 5219
rect 2961 5179 3019 5185
rect 1946 5040 1952 5092
rect 2004 5080 2010 5092
rect 2041 5083 2099 5089
rect 2041 5080 2053 5083
rect 2004 5052 2053 5080
rect 2004 5040 2010 5052
rect 2041 5049 2053 5052
rect 2087 5080 2099 5083
rect 2498 5080 2504 5092
rect 2087 5052 2504 5080
rect 2087 5049 2099 5052
rect 2041 5043 2099 5049
rect 2498 5040 2504 5052
rect 2556 5040 2562 5092
rect 2225 5015 2283 5021
rect 2225 4981 2237 5015
rect 2271 5012 2283 5015
rect 2590 5012 2596 5024
rect 2271 4984 2596 5012
rect 2271 4981 2283 4984
rect 2225 4975 2283 4981
rect 2590 4972 2596 4984
rect 2648 4972 2654 5024
rect 1104 4922 5796 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 5796 4922
rect 1104 4848 5796 4870
rect 4065 4811 4123 4817
rect 4065 4777 4077 4811
rect 4111 4808 4123 4811
rect 4982 4808 4988 4820
rect 4111 4780 4988 4808
rect 4111 4777 4123 4780
rect 4065 4771 4123 4777
rect 4982 4768 4988 4780
rect 5040 4768 5046 4820
rect 14 4700 20 4752
rect 72 4740 78 4752
rect 2409 4743 2467 4749
rect 2409 4740 2421 4743
rect 72 4712 2421 4740
rect 72 4700 78 4712
rect 2409 4709 2421 4712
rect 2455 4709 2467 4743
rect 2409 4703 2467 4709
rect 3050 4632 3056 4684
rect 3108 4672 3114 4684
rect 3108 4644 4016 4672
rect 3108 4632 3114 4644
rect 1854 4564 1860 4616
rect 1912 4564 1918 4616
rect 2590 4564 2596 4616
rect 2648 4604 2654 4616
rect 3068 4604 3096 4632
rect 3988 4616 4016 4644
rect 2648 4576 3096 4604
rect 2648 4564 2654 4576
rect 3142 4564 3148 4616
rect 3200 4564 3206 4616
rect 3970 4564 3976 4616
rect 4028 4564 4034 4616
rect 4706 4564 4712 4616
rect 4764 4604 4770 4616
rect 4801 4607 4859 4613
rect 4801 4604 4813 4607
rect 4764 4576 4813 4604
rect 4764 4564 4770 4576
rect 4801 4573 4813 4576
rect 4847 4573 4859 4607
rect 4801 4567 4859 4573
rect 934 4428 940 4480
rect 992 4468 998 4480
rect 1673 4471 1731 4477
rect 1673 4468 1685 4471
rect 992 4440 1685 4468
rect 992 4428 998 4440
rect 1673 4437 1685 4440
rect 1719 4437 1731 4471
rect 1673 4431 1731 4437
rect 3234 4428 3240 4480
rect 3292 4468 3298 4480
rect 3329 4471 3387 4477
rect 3329 4468 3341 4471
rect 3292 4440 3341 4468
rect 3292 4428 3298 4440
rect 3329 4437 3341 4440
rect 3375 4437 3387 4471
rect 3329 4431 3387 4437
rect 4246 4428 4252 4480
rect 4304 4468 4310 4480
rect 4709 4471 4767 4477
rect 4709 4468 4721 4471
rect 4304 4440 4721 4468
rect 4304 4428 4310 4440
rect 4709 4437 4721 4440
rect 4755 4437 4767 4471
rect 4709 4431 4767 4437
rect 1104 4378 5796 4400
rect 1104 4326 2610 4378
rect 2662 4326 2674 4378
rect 2726 4326 2738 4378
rect 2790 4326 2802 4378
rect 2854 4326 2866 4378
rect 2918 4326 5796 4378
rect 1104 4304 5796 4326
rect 3142 4264 3148 4276
rect 2792 4236 3148 4264
rect 2792 4196 2820 4236
rect 3142 4224 3148 4236
rect 3200 4224 3206 4276
rect 2240 4168 2820 4196
rect 3726 4168 4660 4196
rect 1762 4088 1768 4140
rect 1820 4088 1826 4140
rect 2240 4128 2268 4168
rect 4632 4137 4660 4168
rect 2148 4100 2268 4128
rect 4617 4131 4675 4137
rect 1673 4063 1731 4069
rect 1673 4029 1685 4063
rect 1719 4060 1731 4063
rect 2148 4060 2176 4100
rect 4617 4097 4629 4131
rect 4663 4097 4675 4131
rect 4617 4091 4675 4097
rect 4706 4088 4712 4140
rect 4764 4088 4770 4140
rect 1719 4032 2176 4060
rect 2225 4063 2283 4069
rect 1719 4029 1731 4032
rect 1673 4023 1731 4029
rect 2225 4029 2237 4063
rect 2271 4029 2283 4063
rect 2225 4023 2283 4029
rect 2240 3924 2268 4023
rect 2498 4020 2504 4072
rect 2556 4020 2562 4072
rect 3878 3924 3884 3936
rect 2240 3896 3884 3924
rect 3878 3884 3884 3896
rect 3936 3884 3942 3936
rect 3973 3927 4031 3933
rect 3973 3893 3985 3927
rect 4019 3924 4031 3927
rect 4982 3924 4988 3936
rect 4019 3896 4988 3924
rect 4019 3893 4031 3896
rect 3973 3887 4031 3893
rect 4982 3884 4988 3896
rect 5040 3884 5046 3936
rect 1104 3834 5796 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 5796 3834
rect 1104 3760 5796 3782
rect 1673 3723 1731 3729
rect 1673 3689 1685 3723
rect 1719 3720 1731 3723
rect 1762 3720 1768 3732
rect 1719 3692 1768 3720
rect 1719 3689 1731 3692
rect 1673 3683 1731 3689
rect 1762 3680 1768 3692
rect 1820 3680 1826 3732
rect 2590 3680 2596 3732
rect 2648 3720 2654 3732
rect 2648 3692 5120 3720
rect 2648 3680 2654 3692
rect 3878 3612 3884 3664
rect 3936 3652 3942 3664
rect 3936 3624 4936 3652
rect 3936 3612 3942 3624
rect 4246 3584 4252 3596
rect 2056 3556 4252 3584
rect 2056 3502 2084 3556
rect 4246 3544 4252 3556
rect 4304 3544 4310 3596
rect 3421 3519 3479 3525
rect 3421 3485 3433 3519
rect 3467 3516 3479 3519
rect 3510 3516 3516 3528
rect 3467 3488 3516 3516
rect 3467 3485 3479 3488
rect 3421 3479 3479 3485
rect 3510 3476 3516 3488
rect 3568 3476 3574 3528
rect 4157 3519 4215 3525
rect 4157 3485 4169 3519
rect 4203 3516 4215 3519
rect 4706 3516 4712 3528
rect 4203 3488 4712 3516
rect 4203 3485 4215 3488
rect 4157 3479 4215 3485
rect 4706 3476 4712 3488
rect 4764 3476 4770 3528
rect 4798 3476 4804 3528
rect 4856 3476 4862 3528
rect 3145 3451 3203 3457
rect 3145 3417 3157 3451
rect 3191 3448 3203 3451
rect 4617 3451 4675 3457
rect 4617 3448 4629 3451
rect 3191 3420 4629 3448
rect 3191 3417 3203 3420
rect 3145 3411 3203 3417
rect 4617 3417 4629 3420
rect 4663 3417 4675 3451
rect 4908 3448 4936 3624
rect 5092 3525 5120 3692
rect 5077 3519 5135 3525
rect 5077 3485 5089 3519
rect 5123 3485 5135 3519
rect 5077 3479 5135 3485
rect 5261 3519 5319 3525
rect 5261 3485 5273 3519
rect 5307 3485 5319 3519
rect 5261 3479 5319 3485
rect 5276 3448 5304 3479
rect 4908 3420 5304 3448
rect 4617 3411 4675 3417
rect 1762 3340 1768 3392
rect 1820 3380 1826 3392
rect 3878 3380 3884 3392
rect 1820 3352 3884 3380
rect 1820 3340 1826 3352
rect 3878 3340 3884 3352
rect 3936 3340 3942 3392
rect 4065 3383 4123 3389
rect 4065 3349 4077 3383
rect 4111 3380 4123 3383
rect 4246 3380 4252 3392
rect 4111 3352 4252 3380
rect 4111 3349 4123 3352
rect 4065 3343 4123 3349
rect 4246 3340 4252 3352
rect 4304 3340 4310 3392
rect 1104 3290 5796 3312
rect 1104 3238 2610 3290
rect 2662 3238 2674 3290
rect 2726 3238 2738 3290
rect 2790 3238 2802 3290
rect 2854 3238 2866 3290
rect 2918 3238 5796 3290
rect 1104 3216 5796 3238
rect 3970 3136 3976 3188
rect 4028 3176 4034 3188
rect 5261 3179 5319 3185
rect 5261 3176 5273 3179
rect 4028 3148 5273 3176
rect 4028 3136 4034 3148
rect 5261 3145 5273 3148
rect 5307 3145 5319 3179
rect 5261 3139 5319 3145
rect 3786 3068 3792 3120
rect 3844 3068 3850 3120
rect 4246 3068 4252 3120
rect 4304 3068 4310 3120
rect 2225 3043 2283 3049
rect 2225 3009 2237 3043
rect 2271 3040 2283 3043
rect 2406 3040 2412 3052
rect 2271 3012 2412 3040
rect 2271 3009 2283 3012
rect 2225 3003 2283 3009
rect 2406 3000 2412 3012
rect 2464 3000 2470 3052
rect 2314 2932 2320 2984
rect 2372 2972 2378 2984
rect 2372 2944 2452 2972
rect 2372 2932 2378 2944
rect 2424 2836 2452 2944
rect 2498 2932 2504 2984
rect 2556 2972 2562 2984
rect 2593 2975 2651 2981
rect 2593 2972 2605 2975
rect 2556 2944 2605 2972
rect 2556 2932 2562 2944
rect 2593 2941 2605 2944
rect 2639 2941 2651 2975
rect 2593 2935 2651 2941
rect 3510 2932 3516 2984
rect 3568 2932 3574 2984
rect 4982 2836 4988 2848
rect 2424 2808 4988 2836
rect 4982 2796 4988 2808
rect 5040 2796 5046 2848
rect 1104 2746 5796 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 5796 2746
rect 1104 2672 5796 2694
rect 2133 2635 2191 2641
rect 2133 2601 2145 2635
rect 2179 2632 2191 2635
rect 3510 2632 3516 2644
rect 2179 2604 3516 2632
rect 2179 2601 2191 2604
rect 2133 2595 2191 2601
rect 3510 2592 3516 2604
rect 3568 2592 3574 2644
rect 5169 2635 5227 2641
rect 5169 2601 5181 2635
rect 5215 2632 5227 2635
rect 5442 2632 5448 2644
rect 5215 2604 5448 2632
rect 5215 2601 5227 2604
rect 5169 2595 5227 2601
rect 5442 2592 5448 2604
rect 5500 2592 5506 2644
rect 3421 2431 3479 2437
rect 3421 2397 3433 2431
rect 3467 2428 3479 2431
rect 4062 2428 4068 2440
rect 3467 2400 4068 2428
rect 3467 2397 3479 2400
rect 3421 2391 3479 2397
rect 4062 2388 4068 2400
rect 4120 2388 4126 2440
rect 4522 2388 4528 2440
rect 4580 2388 4586 2440
rect 4982 2388 4988 2440
rect 5040 2388 5046 2440
rect 4341 2295 4399 2301
rect 4341 2261 4353 2295
rect 4387 2292 4399 2295
rect 6454 2292 6460 2304
rect 4387 2264 6460 2292
rect 4387 2261 4399 2264
rect 4341 2255 4399 2261
rect 6454 2252 6460 2264
rect 6512 2252 6518 2304
rect 1104 2202 5796 2224
rect 1104 2150 2610 2202
rect 2662 2150 2674 2202
rect 2726 2150 2738 2202
rect 2790 2150 2802 2202
rect 2854 2150 2866 2202
rect 2918 2150 5796 2202
rect 1104 2128 5796 2150
<< via1 >>
rect 1950 9222 2002 9274
rect 2014 9222 2066 9274
rect 2078 9222 2130 9274
rect 2142 9222 2194 9274
rect 2206 9222 2258 9274
rect 5172 9163 5224 9172
rect 5172 9129 5181 9163
rect 5181 9129 5215 9163
rect 5215 9129 5224 9163
rect 5172 9120 5224 9129
rect 2964 9052 3016 9104
rect 1860 8984 1912 9036
rect 2412 8916 2464 8968
rect 4252 8959 4304 8968
rect 4252 8925 4261 8959
rect 4261 8925 4295 8959
rect 4295 8925 4304 8959
rect 4252 8916 4304 8925
rect 4344 8916 4396 8968
rect 3056 8848 3108 8900
rect 2610 8678 2662 8730
rect 2674 8678 2726 8730
rect 2738 8678 2790 8730
rect 2802 8678 2854 8730
rect 2866 8678 2918 8730
rect 940 8576 992 8628
rect 5908 8576 5960 8628
rect 2504 8440 2556 8492
rect 4988 8483 5040 8492
rect 4988 8449 4997 8483
rect 4997 8449 5031 8483
rect 5031 8449 5040 8483
rect 4988 8440 5040 8449
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 2610 7590 2662 7642
rect 2674 7590 2726 7642
rect 2738 7590 2790 7642
rect 2802 7590 2854 7642
rect 2866 7590 2918 7642
rect 4896 7352 4948 7404
rect 3792 7327 3844 7336
rect 3792 7293 3801 7327
rect 3801 7293 3835 7327
rect 3835 7293 3844 7327
rect 3792 7284 3844 7293
rect 3884 7148 3936 7200
rect 5264 7191 5316 7200
rect 5264 7157 5273 7191
rect 5273 7157 5307 7191
rect 5307 7157 5316 7191
rect 5264 7148 5316 7157
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 1768 6808 1820 6860
rect 4344 6808 4396 6860
rect 4896 6851 4948 6860
rect 4896 6817 4905 6851
rect 4905 6817 4939 6851
rect 4939 6817 4948 6851
rect 4896 6808 4948 6817
rect 2228 6740 2280 6792
rect 4252 6740 4304 6792
rect 4712 6740 4764 6792
rect 3056 6672 3108 6724
rect 2412 6604 2464 6656
rect 4160 6604 4212 6656
rect 2610 6502 2662 6554
rect 2674 6502 2726 6554
rect 2738 6502 2790 6554
rect 2802 6502 2854 6554
rect 2866 6502 2918 6554
rect 2320 6264 2372 6316
rect 4068 6264 4120 6316
rect 5908 6264 5960 6316
rect 4712 6128 4764 6180
rect 1860 6060 1912 6112
rect 3884 6103 3936 6112
rect 3884 6069 3893 6103
rect 3893 6069 3927 6103
rect 3927 6069 3936 6103
rect 3884 6060 3936 6069
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 3792 5788 3844 5840
rect 2504 5720 2556 5772
rect 1952 5652 2004 5704
rect 2872 5652 2924 5704
rect 4160 5720 4212 5772
rect 4804 5720 4856 5772
rect 4528 5652 4580 5704
rect 5264 5652 5316 5704
rect 3792 5516 3844 5568
rect 2610 5414 2662 5466
rect 2674 5414 2726 5466
rect 2738 5414 2790 5466
rect 2802 5414 2854 5466
rect 2866 5414 2918 5466
rect 4068 5312 4120 5364
rect 2320 5244 2372 5296
rect 2412 5287 2464 5296
rect 2412 5253 2421 5287
rect 2421 5253 2455 5287
rect 2455 5253 2464 5287
rect 2412 5244 2464 5253
rect 940 5176 992 5228
rect 1952 5040 2004 5092
rect 2504 5040 2556 5092
rect 2596 4972 2648 5024
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 4988 4768 5040 4820
rect 20 4700 72 4752
rect 3056 4632 3108 4684
rect 1860 4607 1912 4616
rect 1860 4573 1869 4607
rect 1869 4573 1903 4607
rect 1903 4573 1912 4607
rect 1860 4564 1912 4573
rect 2596 4607 2648 4616
rect 2596 4573 2605 4607
rect 2605 4573 2639 4607
rect 2639 4573 2648 4607
rect 2596 4564 2648 4573
rect 3148 4607 3200 4616
rect 3148 4573 3157 4607
rect 3157 4573 3191 4607
rect 3191 4573 3200 4607
rect 3148 4564 3200 4573
rect 3976 4607 4028 4616
rect 3976 4573 3985 4607
rect 3985 4573 4019 4607
rect 4019 4573 4028 4607
rect 3976 4564 4028 4573
rect 4712 4564 4764 4616
rect 940 4428 992 4480
rect 3240 4428 3292 4480
rect 4252 4428 4304 4480
rect 2610 4326 2662 4378
rect 2674 4326 2726 4378
rect 2738 4326 2790 4378
rect 2802 4326 2854 4378
rect 2866 4326 2918 4378
rect 3148 4224 3200 4276
rect 1768 4131 1820 4140
rect 1768 4097 1777 4131
rect 1777 4097 1811 4131
rect 1811 4097 1820 4131
rect 1768 4088 1820 4097
rect 4712 4131 4764 4140
rect 4712 4097 4721 4131
rect 4721 4097 4755 4131
rect 4755 4097 4764 4131
rect 4712 4088 4764 4097
rect 2504 4063 2556 4072
rect 2504 4029 2513 4063
rect 2513 4029 2547 4063
rect 2547 4029 2556 4063
rect 2504 4020 2556 4029
rect 3884 3884 3936 3936
rect 4988 3884 5040 3936
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 1768 3680 1820 3732
rect 2596 3680 2648 3732
rect 3884 3612 3936 3664
rect 4252 3544 4304 3596
rect 3516 3476 3568 3528
rect 4712 3476 4764 3528
rect 4804 3519 4856 3528
rect 4804 3485 4813 3519
rect 4813 3485 4847 3519
rect 4847 3485 4856 3519
rect 4804 3476 4856 3485
rect 1768 3340 1820 3392
rect 3884 3340 3936 3392
rect 4252 3340 4304 3392
rect 2610 3238 2662 3290
rect 2674 3238 2726 3290
rect 2738 3238 2790 3290
rect 2802 3238 2854 3290
rect 2866 3238 2918 3290
rect 3976 3136 4028 3188
rect 3792 3111 3844 3120
rect 3792 3077 3801 3111
rect 3801 3077 3835 3111
rect 3835 3077 3844 3111
rect 3792 3068 3844 3077
rect 4252 3068 4304 3120
rect 2412 3000 2464 3052
rect 2320 2975 2372 2984
rect 2320 2941 2329 2975
rect 2329 2941 2363 2975
rect 2363 2941 2372 2975
rect 2320 2932 2372 2941
rect 2504 2932 2556 2984
rect 3516 2975 3568 2984
rect 3516 2941 3525 2975
rect 3525 2941 3559 2975
rect 3559 2941 3568 2975
rect 3516 2932 3568 2941
rect 4988 2796 5040 2848
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 3516 2592 3568 2644
rect 5448 2592 5500 2644
rect 4068 2388 4120 2440
rect 4528 2431 4580 2440
rect 4528 2397 4537 2431
rect 4537 2397 4571 2431
rect 4571 2397 4580 2431
rect 4528 2388 4580 2397
rect 4988 2431 5040 2440
rect 4988 2397 4997 2431
rect 4997 2397 5031 2431
rect 5031 2397 5040 2431
rect 4988 2388 5040 2397
rect 6460 2252 6512 2304
rect 2610 2150 2662 2202
rect 2674 2150 2726 2202
rect 2738 2150 2790 2202
rect 2802 2150 2854 2202
rect 2866 2150 2918 2202
<< metal2 >>
rect 1950 10624 2006 11424
rect 5170 10624 5226 11424
rect 938 10296 994 10305
rect 938 10231 994 10240
rect 952 8634 980 10231
rect 1964 9466 1992 10624
rect 1872 9438 1992 9466
rect 1872 9042 1900 9438
rect 1950 9276 2258 9285
rect 1950 9274 1956 9276
rect 2012 9274 2036 9276
rect 2092 9274 2116 9276
rect 2172 9274 2196 9276
rect 2252 9274 2258 9276
rect 2012 9222 2014 9274
rect 2194 9222 2196 9274
rect 1950 9220 1956 9222
rect 2012 9220 2036 9222
rect 2092 9220 2116 9222
rect 2172 9220 2196 9222
rect 2252 9220 2258 9222
rect 1950 9211 2258 9220
rect 5184 9178 5212 10624
rect 5906 9616 5962 9625
rect 5906 9551 5962 9560
rect 5172 9172 5224 9178
rect 5172 9114 5224 9120
rect 2964 9104 3016 9110
rect 2964 9046 3016 9052
rect 1860 9036 1912 9042
rect 1860 8978 1912 8984
rect 2412 8968 2464 8974
rect 2412 8910 2464 8916
rect 940 8628 992 8634
rect 940 8570 992 8576
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 938 6896 994 6905
rect 938 6831 994 6840
rect 1768 6860 1820 6866
rect 952 5234 980 6831
rect 1768 6802 1820 6808
rect 940 5228 992 5234
rect 940 5170 992 5176
rect 20 4752 72 4758
rect 20 4694 72 4700
rect 32 800 60 4694
rect 940 4480 992 4486
rect 940 4422 992 4428
rect 952 3505 980 4422
rect 1780 4146 1808 6802
rect 2228 6792 2280 6798
rect 2280 6740 2360 6746
rect 2228 6734 2360 6740
rect 2240 6718 2360 6734
rect 2332 6322 2360 6718
rect 2424 6662 2452 8910
rect 2610 8732 2918 8741
rect 2610 8730 2616 8732
rect 2672 8730 2696 8732
rect 2752 8730 2776 8732
rect 2832 8730 2856 8732
rect 2912 8730 2918 8732
rect 2672 8678 2674 8730
rect 2854 8678 2856 8730
rect 2610 8676 2616 8678
rect 2672 8676 2696 8678
rect 2752 8676 2776 8678
rect 2832 8676 2856 8678
rect 2912 8676 2918 8678
rect 2610 8667 2918 8676
rect 2504 8492 2556 8498
rect 2504 8434 2556 8440
rect 2412 6656 2464 6662
rect 2412 6598 2464 6604
rect 2320 6316 2372 6322
rect 2320 6258 2372 6264
rect 1860 6112 1912 6118
rect 1860 6054 1912 6060
rect 1872 4622 1900 6054
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 1952 5704 2004 5710
rect 1952 5646 2004 5652
rect 1964 5098 1992 5646
rect 2332 5302 2360 6258
rect 2424 5302 2452 6598
rect 2516 5778 2544 8434
rect 2610 7644 2918 7653
rect 2610 7642 2616 7644
rect 2672 7642 2696 7644
rect 2752 7642 2776 7644
rect 2832 7642 2856 7644
rect 2912 7642 2918 7644
rect 2672 7590 2674 7642
rect 2854 7590 2856 7642
rect 2610 7588 2616 7590
rect 2672 7588 2696 7590
rect 2752 7588 2776 7590
rect 2832 7588 2856 7590
rect 2912 7588 2918 7590
rect 2610 7579 2918 7588
rect 2610 6556 2918 6565
rect 2610 6554 2616 6556
rect 2672 6554 2696 6556
rect 2752 6554 2776 6556
rect 2832 6554 2856 6556
rect 2912 6554 2918 6556
rect 2672 6502 2674 6554
rect 2854 6502 2856 6554
rect 2610 6500 2616 6502
rect 2672 6500 2696 6502
rect 2752 6500 2776 6502
rect 2832 6500 2856 6502
rect 2912 6500 2918 6502
rect 2610 6491 2918 6500
rect 2976 6338 3004 9046
rect 4252 8968 4304 8974
rect 4252 8910 4304 8916
rect 4344 8968 4396 8974
rect 4344 8910 4396 8916
rect 3056 8900 3108 8906
rect 3056 8842 3108 8848
rect 3068 6730 3096 8842
rect 3792 7336 3844 7342
rect 3792 7278 3844 7284
rect 3056 6724 3108 6730
rect 3056 6666 3108 6672
rect 2884 6310 3004 6338
rect 2504 5772 2556 5778
rect 2504 5714 2556 5720
rect 2884 5710 2912 6310
rect 2872 5704 2924 5710
rect 2872 5646 2924 5652
rect 2610 5468 2918 5477
rect 2610 5466 2616 5468
rect 2672 5466 2696 5468
rect 2752 5466 2776 5468
rect 2832 5466 2856 5468
rect 2912 5466 2918 5468
rect 2672 5414 2674 5466
rect 2854 5414 2856 5466
rect 2610 5412 2616 5414
rect 2672 5412 2696 5414
rect 2752 5412 2776 5414
rect 2832 5412 2856 5414
rect 2912 5412 2918 5414
rect 2610 5403 2918 5412
rect 2320 5296 2372 5302
rect 2320 5238 2372 5244
rect 2412 5296 2464 5302
rect 2412 5238 2464 5244
rect 1952 5092 2004 5098
rect 1952 5034 2004 5040
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 1860 4616 1912 4622
rect 1860 4558 1912 4564
rect 1768 4140 1820 4146
rect 1768 4082 1820 4088
rect 1780 3738 1808 4082
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 1768 3732 1820 3738
rect 1768 3674 1820 3680
rect 938 3496 994 3505
rect 938 3431 994 3440
rect 1780 3398 1808 3674
rect 1768 3392 1820 3398
rect 1768 3334 1820 3340
rect 2332 2990 2360 5238
rect 2424 3058 2452 5238
rect 2504 5092 2556 5098
rect 2504 5034 2556 5040
rect 2516 4162 2544 5034
rect 2596 5024 2648 5030
rect 2596 4966 2648 4972
rect 2608 4622 2636 4966
rect 3068 4690 3096 6666
rect 3804 5846 3832 7278
rect 3884 7200 3936 7206
rect 3884 7142 3936 7148
rect 3896 6118 3924 7142
rect 4264 6798 4292 8910
rect 4356 6866 4384 8910
rect 5920 8634 5948 9551
rect 5908 8628 5960 8634
rect 5908 8570 5960 8576
rect 4988 8492 5040 8498
rect 4988 8434 5040 8440
rect 4896 7404 4948 7410
rect 4896 7346 4948 7352
rect 4908 6866 4936 7346
rect 4344 6860 4396 6866
rect 4344 6802 4396 6808
rect 4896 6860 4948 6866
rect 4896 6802 4948 6808
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 4712 6792 4764 6798
rect 4712 6734 4764 6740
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 4068 6316 4120 6322
rect 4068 6258 4120 6264
rect 3884 6112 3936 6118
rect 3884 6054 3936 6060
rect 3792 5840 3844 5846
rect 3792 5782 3844 5788
rect 3792 5568 3844 5574
rect 3792 5510 3844 5516
rect 3056 4684 3108 4690
rect 3056 4626 3108 4632
rect 2596 4616 2648 4622
rect 2596 4558 2648 4564
rect 3148 4616 3200 4622
rect 3148 4558 3200 4564
rect 2610 4380 2918 4389
rect 2610 4378 2616 4380
rect 2672 4378 2696 4380
rect 2752 4378 2776 4380
rect 2832 4378 2856 4380
rect 2912 4378 2918 4380
rect 2672 4326 2674 4378
rect 2854 4326 2856 4378
rect 2610 4324 2616 4326
rect 2672 4324 2696 4326
rect 2752 4324 2776 4326
rect 2832 4324 2856 4326
rect 2912 4324 2918 4326
rect 2610 4315 2918 4324
rect 3160 4282 3188 4558
rect 3240 4480 3292 4486
rect 3240 4422 3292 4428
rect 3148 4276 3200 4282
rect 3148 4218 3200 4224
rect 2516 4134 2636 4162
rect 2504 4072 2556 4078
rect 2504 4014 2556 4020
rect 2412 3052 2464 3058
rect 2412 2994 2464 3000
rect 2516 2990 2544 4014
rect 2608 3738 2636 4134
rect 2596 3732 2648 3738
rect 2596 3674 2648 3680
rect 2610 3292 2918 3301
rect 2610 3290 2616 3292
rect 2672 3290 2696 3292
rect 2752 3290 2776 3292
rect 2832 3290 2856 3292
rect 2912 3290 2918 3292
rect 2672 3238 2674 3290
rect 2854 3238 2856 3290
rect 2610 3236 2616 3238
rect 2672 3236 2696 3238
rect 2752 3236 2776 3238
rect 2832 3236 2856 3238
rect 2912 3236 2918 3238
rect 2610 3227 2918 3236
rect 2320 2984 2372 2990
rect 2320 2926 2372 2932
rect 2504 2984 2556 2990
rect 2504 2926 2556 2932
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 2610 2204 2918 2213
rect 2610 2202 2616 2204
rect 2672 2202 2696 2204
rect 2752 2202 2776 2204
rect 2832 2202 2856 2204
rect 2912 2202 2918 2204
rect 2672 2150 2674 2202
rect 2854 2150 2856 2202
rect 2610 2148 2616 2150
rect 2672 2148 2696 2150
rect 2752 2148 2776 2150
rect 2832 2148 2856 2150
rect 2912 2148 2918 2150
rect 2610 2139 2918 2148
rect 3252 800 3280 4422
rect 3516 3528 3568 3534
rect 3516 3470 3568 3476
rect 3528 2990 3556 3470
rect 3804 3126 3832 5510
rect 3896 3942 3924 6054
rect 4080 5370 4108 6258
rect 4172 5778 4200 6598
rect 4724 6186 4752 6734
rect 4712 6180 4764 6186
rect 4712 6122 4764 6128
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 4528 5704 4580 5710
rect 4528 5646 4580 5652
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 3884 3936 3936 3942
rect 3884 3878 3936 3884
rect 3884 3664 3936 3670
rect 3884 3606 3936 3612
rect 3896 3398 3924 3606
rect 3884 3392 3936 3398
rect 3884 3334 3936 3340
rect 3988 3194 4016 4558
rect 3976 3188 4028 3194
rect 3976 3130 4028 3136
rect 3792 3120 3844 3126
rect 3792 3062 3844 3068
rect 3516 2984 3568 2990
rect 3516 2926 3568 2932
rect 3528 2650 3556 2926
rect 3516 2644 3568 2650
rect 3516 2586 3568 2592
rect 4080 2446 4108 5306
rect 4252 4480 4304 4486
rect 4252 4422 4304 4428
rect 4264 3602 4292 4422
rect 4252 3596 4304 3602
rect 4252 3538 4304 3544
rect 4252 3392 4304 3398
rect 4252 3334 4304 3340
rect 4264 3126 4292 3334
rect 4252 3120 4304 3126
rect 4252 3062 4304 3068
rect 4540 2446 4568 5646
rect 4724 4622 4752 6122
rect 4804 5772 4856 5778
rect 4804 5714 4856 5720
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 4724 4146 4752 4558
rect 4712 4140 4764 4146
rect 4712 4082 4764 4088
rect 4724 3534 4752 4082
rect 4816 3534 4844 5714
rect 5000 4826 5028 8434
rect 5264 7200 5316 7206
rect 5264 7142 5316 7148
rect 5276 5710 5304 7142
rect 5908 6316 5960 6322
rect 5908 6258 5960 6264
rect 5920 6225 5948 6258
rect 5906 6216 5962 6225
rect 5906 6151 5962 6160
rect 5264 5704 5316 5710
rect 5264 5646 5316 5652
rect 4988 4820 5040 4826
rect 4988 4762 5040 4768
rect 4988 3936 5040 3942
rect 4988 3878 5040 3884
rect 4712 3528 4764 3534
rect 4712 3470 4764 3476
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 5000 2854 5028 3878
rect 4988 2848 5040 2854
rect 4988 2790 5040 2796
rect 5446 2816 5502 2825
rect 5000 2446 5028 2790
rect 5446 2751 5502 2760
rect 5460 2650 5488 2751
rect 5448 2644 5500 2650
rect 5448 2586 5500 2592
rect 4068 2440 4120 2446
rect 4068 2382 4120 2388
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 4988 2440 5040 2446
rect 4988 2382 5040 2388
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 6472 800 6500 2246
rect 18 0 74 800
rect 3238 0 3294 800
rect 6458 0 6514 800
<< via2 >>
rect 938 10240 994 10296
rect 1956 9274 2012 9276
rect 2036 9274 2092 9276
rect 2116 9274 2172 9276
rect 2196 9274 2252 9276
rect 1956 9222 2002 9274
rect 2002 9222 2012 9274
rect 2036 9222 2066 9274
rect 2066 9222 2078 9274
rect 2078 9222 2092 9274
rect 2116 9222 2130 9274
rect 2130 9222 2142 9274
rect 2142 9222 2172 9274
rect 2196 9222 2206 9274
rect 2206 9222 2252 9274
rect 1956 9220 2012 9222
rect 2036 9220 2092 9222
rect 2116 9220 2172 9222
rect 2196 9220 2252 9222
rect 5906 9560 5962 9616
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 938 6840 994 6896
rect 2616 8730 2672 8732
rect 2696 8730 2752 8732
rect 2776 8730 2832 8732
rect 2856 8730 2912 8732
rect 2616 8678 2662 8730
rect 2662 8678 2672 8730
rect 2696 8678 2726 8730
rect 2726 8678 2738 8730
rect 2738 8678 2752 8730
rect 2776 8678 2790 8730
rect 2790 8678 2802 8730
rect 2802 8678 2832 8730
rect 2856 8678 2866 8730
rect 2866 8678 2912 8730
rect 2616 8676 2672 8678
rect 2696 8676 2752 8678
rect 2776 8676 2832 8678
rect 2856 8676 2912 8678
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 2616 7642 2672 7644
rect 2696 7642 2752 7644
rect 2776 7642 2832 7644
rect 2856 7642 2912 7644
rect 2616 7590 2662 7642
rect 2662 7590 2672 7642
rect 2696 7590 2726 7642
rect 2726 7590 2738 7642
rect 2738 7590 2752 7642
rect 2776 7590 2790 7642
rect 2790 7590 2802 7642
rect 2802 7590 2832 7642
rect 2856 7590 2866 7642
rect 2866 7590 2912 7642
rect 2616 7588 2672 7590
rect 2696 7588 2752 7590
rect 2776 7588 2832 7590
rect 2856 7588 2912 7590
rect 2616 6554 2672 6556
rect 2696 6554 2752 6556
rect 2776 6554 2832 6556
rect 2856 6554 2912 6556
rect 2616 6502 2662 6554
rect 2662 6502 2672 6554
rect 2696 6502 2726 6554
rect 2726 6502 2738 6554
rect 2738 6502 2752 6554
rect 2776 6502 2790 6554
rect 2790 6502 2802 6554
rect 2802 6502 2832 6554
rect 2856 6502 2866 6554
rect 2866 6502 2912 6554
rect 2616 6500 2672 6502
rect 2696 6500 2752 6502
rect 2776 6500 2832 6502
rect 2856 6500 2912 6502
rect 2616 5466 2672 5468
rect 2696 5466 2752 5468
rect 2776 5466 2832 5468
rect 2856 5466 2912 5468
rect 2616 5414 2662 5466
rect 2662 5414 2672 5466
rect 2696 5414 2726 5466
rect 2726 5414 2738 5466
rect 2738 5414 2752 5466
rect 2776 5414 2790 5466
rect 2790 5414 2802 5466
rect 2802 5414 2832 5466
rect 2856 5414 2866 5466
rect 2866 5414 2912 5466
rect 2616 5412 2672 5414
rect 2696 5412 2752 5414
rect 2776 5412 2832 5414
rect 2856 5412 2912 5414
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 938 3440 994 3496
rect 2616 4378 2672 4380
rect 2696 4378 2752 4380
rect 2776 4378 2832 4380
rect 2856 4378 2912 4380
rect 2616 4326 2662 4378
rect 2662 4326 2672 4378
rect 2696 4326 2726 4378
rect 2726 4326 2738 4378
rect 2738 4326 2752 4378
rect 2776 4326 2790 4378
rect 2790 4326 2802 4378
rect 2802 4326 2832 4378
rect 2856 4326 2866 4378
rect 2866 4326 2912 4378
rect 2616 4324 2672 4326
rect 2696 4324 2752 4326
rect 2776 4324 2832 4326
rect 2856 4324 2912 4326
rect 2616 3290 2672 3292
rect 2696 3290 2752 3292
rect 2776 3290 2832 3292
rect 2856 3290 2912 3292
rect 2616 3238 2662 3290
rect 2662 3238 2672 3290
rect 2696 3238 2726 3290
rect 2726 3238 2738 3290
rect 2738 3238 2752 3290
rect 2776 3238 2790 3290
rect 2790 3238 2802 3290
rect 2802 3238 2832 3290
rect 2856 3238 2866 3290
rect 2866 3238 2912 3290
rect 2616 3236 2672 3238
rect 2696 3236 2752 3238
rect 2776 3236 2832 3238
rect 2856 3236 2912 3238
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 2616 2202 2672 2204
rect 2696 2202 2752 2204
rect 2776 2202 2832 2204
rect 2856 2202 2912 2204
rect 2616 2150 2662 2202
rect 2662 2150 2672 2202
rect 2696 2150 2726 2202
rect 2726 2150 2738 2202
rect 2738 2150 2752 2202
rect 2776 2150 2790 2202
rect 2790 2150 2802 2202
rect 2802 2150 2832 2202
rect 2856 2150 2866 2202
rect 2866 2150 2912 2202
rect 2616 2148 2672 2150
rect 2696 2148 2752 2150
rect 2776 2148 2832 2150
rect 2856 2148 2912 2150
rect 5906 6160 5962 6216
rect 5446 2760 5502 2816
<< metal3 >>
rect 0 10298 800 10328
rect 933 10298 999 10301
rect 0 10296 999 10298
rect 0 10240 938 10296
rect 994 10240 999 10296
rect 0 10238 999 10240
rect 0 10208 800 10238
rect 933 10235 999 10238
rect 5901 9618 5967 9621
rect 6100 9618 6900 9648
rect 5901 9616 6900 9618
rect 5901 9560 5906 9616
rect 5962 9560 6900 9616
rect 5901 9558 6900 9560
rect 5901 9555 5967 9558
rect 6100 9528 6900 9558
rect 1946 9280 2262 9281
rect 1946 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2262 9280
rect 1946 9215 2262 9216
rect 2606 8736 2922 8737
rect 2606 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2922 8736
rect 2606 8671 2922 8672
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 2606 7648 2922 7649
rect 2606 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2922 7648
rect 2606 7583 2922 7584
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 0 6898 800 6928
rect 933 6898 999 6901
rect 0 6896 999 6898
rect 0 6840 938 6896
rect 994 6840 999 6896
rect 0 6838 999 6840
rect 0 6808 800 6838
rect 933 6835 999 6838
rect 2606 6560 2922 6561
rect 2606 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2922 6560
rect 2606 6495 2922 6496
rect 5901 6218 5967 6221
rect 6100 6218 6900 6248
rect 5901 6216 6900 6218
rect 5901 6160 5906 6216
rect 5962 6160 6900 6216
rect 5901 6158 6900 6160
rect 5901 6155 5967 6158
rect 6100 6128 6900 6158
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 2606 5472 2922 5473
rect 2606 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2922 5472
rect 2606 5407 2922 5408
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 2606 4384 2922 4385
rect 2606 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2922 4384
rect 2606 4319 2922 4320
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 0 3498 800 3528
rect 933 3498 999 3501
rect 0 3496 999 3498
rect 0 3440 938 3496
rect 994 3440 999 3496
rect 0 3438 999 3440
rect 0 3408 800 3438
rect 933 3435 999 3438
rect 2606 3296 2922 3297
rect 2606 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2922 3296
rect 2606 3231 2922 3232
rect 5441 2818 5507 2821
rect 6100 2818 6900 2848
rect 5441 2816 6900 2818
rect 5441 2760 5446 2816
rect 5502 2760 6900 2816
rect 5441 2758 6900 2760
rect 5441 2755 5507 2758
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 6100 2728 6900 2758
rect 1946 2687 2262 2688
rect 2606 2208 2922 2209
rect 2606 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2922 2208
rect 2606 2143 2922 2144
<< via3 >>
rect 1952 9276 2016 9280
rect 1952 9220 1956 9276
rect 1956 9220 2012 9276
rect 2012 9220 2016 9276
rect 1952 9216 2016 9220
rect 2032 9276 2096 9280
rect 2032 9220 2036 9276
rect 2036 9220 2092 9276
rect 2092 9220 2096 9276
rect 2032 9216 2096 9220
rect 2112 9276 2176 9280
rect 2112 9220 2116 9276
rect 2116 9220 2172 9276
rect 2172 9220 2176 9276
rect 2112 9216 2176 9220
rect 2192 9276 2256 9280
rect 2192 9220 2196 9276
rect 2196 9220 2252 9276
rect 2252 9220 2256 9276
rect 2192 9216 2256 9220
rect 2612 8732 2676 8736
rect 2612 8676 2616 8732
rect 2616 8676 2672 8732
rect 2672 8676 2676 8732
rect 2612 8672 2676 8676
rect 2692 8732 2756 8736
rect 2692 8676 2696 8732
rect 2696 8676 2752 8732
rect 2752 8676 2756 8732
rect 2692 8672 2756 8676
rect 2772 8732 2836 8736
rect 2772 8676 2776 8732
rect 2776 8676 2832 8732
rect 2832 8676 2836 8732
rect 2772 8672 2836 8676
rect 2852 8732 2916 8736
rect 2852 8676 2856 8732
rect 2856 8676 2912 8732
rect 2912 8676 2916 8732
rect 2852 8672 2916 8676
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 2612 7644 2676 7648
rect 2612 7588 2616 7644
rect 2616 7588 2672 7644
rect 2672 7588 2676 7644
rect 2612 7584 2676 7588
rect 2692 7644 2756 7648
rect 2692 7588 2696 7644
rect 2696 7588 2752 7644
rect 2752 7588 2756 7644
rect 2692 7584 2756 7588
rect 2772 7644 2836 7648
rect 2772 7588 2776 7644
rect 2776 7588 2832 7644
rect 2832 7588 2836 7644
rect 2772 7584 2836 7588
rect 2852 7644 2916 7648
rect 2852 7588 2856 7644
rect 2856 7588 2912 7644
rect 2912 7588 2916 7644
rect 2852 7584 2916 7588
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 2612 6556 2676 6560
rect 2612 6500 2616 6556
rect 2616 6500 2672 6556
rect 2672 6500 2676 6556
rect 2612 6496 2676 6500
rect 2692 6556 2756 6560
rect 2692 6500 2696 6556
rect 2696 6500 2752 6556
rect 2752 6500 2756 6556
rect 2692 6496 2756 6500
rect 2772 6556 2836 6560
rect 2772 6500 2776 6556
rect 2776 6500 2832 6556
rect 2832 6500 2836 6556
rect 2772 6496 2836 6500
rect 2852 6556 2916 6560
rect 2852 6500 2856 6556
rect 2856 6500 2912 6556
rect 2912 6500 2916 6556
rect 2852 6496 2916 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 2612 5468 2676 5472
rect 2612 5412 2616 5468
rect 2616 5412 2672 5468
rect 2672 5412 2676 5468
rect 2612 5408 2676 5412
rect 2692 5468 2756 5472
rect 2692 5412 2696 5468
rect 2696 5412 2752 5468
rect 2752 5412 2756 5468
rect 2692 5408 2756 5412
rect 2772 5468 2836 5472
rect 2772 5412 2776 5468
rect 2776 5412 2832 5468
rect 2832 5412 2836 5468
rect 2772 5408 2836 5412
rect 2852 5468 2916 5472
rect 2852 5412 2856 5468
rect 2856 5412 2912 5468
rect 2912 5412 2916 5468
rect 2852 5408 2916 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 2612 4380 2676 4384
rect 2612 4324 2616 4380
rect 2616 4324 2672 4380
rect 2672 4324 2676 4380
rect 2612 4320 2676 4324
rect 2692 4380 2756 4384
rect 2692 4324 2696 4380
rect 2696 4324 2752 4380
rect 2752 4324 2756 4380
rect 2692 4320 2756 4324
rect 2772 4380 2836 4384
rect 2772 4324 2776 4380
rect 2776 4324 2832 4380
rect 2832 4324 2836 4380
rect 2772 4320 2836 4324
rect 2852 4380 2916 4384
rect 2852 4324 2856 4380
rect 2856 4324 2912 4380
rect 2912 4324 2916 4380
rect 2852 4320 2916 4324
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 2612 3292 2676 3296
rect 2612 3236 2616 3292
rect 2616 3236 2672 3292
rect 2672 3236 2676 3292
rect 2612 3232 2676 3236
rect 2692 3292 2756 3296
rect 2692 3236 2696 3292
rect 2696 3236 2752 3292
rect 2752 3236 2756 3292
rect 2692 3232 2756 3236
rect 2772 3292 2836 3296
rect 2772 3236 2776 3292
rect 2776 3236 2832 3292
rect 2832 3236 2836 3292
rect 2772 3232 2836 3236
rect 2852 3292 2916 3296
rect 2852 3236 2856 3292
rect 2856 3236 2912 3292
rect 2912 3236 2916 3292
rect 2852 3232 2916 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 2612 2204 2676 2208
rect 2612 2148 2616 2204
rect 2616 2148 2672 2204
rect 2672 2148 2676 2204
rect 2612 2144 2676 2148
rect 2692 2204 2756 2208
rect 2692 2148 2696 2204
rect 2696 2148 2752 2204
rect 2752 2148 2756 2204
rect 2692 2144 2756 2148
rect 2772 2204 2836 2208
rect 2772 2148 2776 2204
rect 2776 2148 2832 2204
rect 2832 2148 2836 2204
rect 2772 2144 2836 2148
rect 2852 2204 2916 2208
rect 2852 2148 2856 2204
rect 2856 2148 2912 2204
rect 2912 2148 2916 2204
rect 2852 2144 2916 2148
<< metal4 >>
rect 1944 9280 2264 9296
rect 1944 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2264 9280
rect 1944 8192 2264 9216
rect 1944 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2264 8192
rect 1944 7104 2264 8128
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 2752 2264 3776
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 2128 2264 2688
rect 2604 8736 2924 9296
rect 2604 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2924 8736
rect 2604 7648 2924 8672
rect 2604 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2924 7648
rect 2604 6560 2924 7584
rect 2604 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2924 6560
rect 2604 5472 2924 6496
rect 2604 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2924 5472
rect 2604 4384 2924 5408
rect 2604 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2924 4384
rect 2604 3296 2924 4320
rect 2604 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2924 3296
rect 2604 2208 2924 3232
rect 2604 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2924 2208
rect 2604 2128 2924 2144
use sky130_fd_sc_hd__decap_3  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4140 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38
timestamp 1676037725
transform 1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46
timestamp 1676037725
transform 1 0 5336 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_9
timestamp 1676037725
transform 1 0 1932 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_17 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2668 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_25
timestamp 1676037725
transform 1 0 3404 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_46
timestamp 1676037725
transform 1 0 5336 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1676037725
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_34
timestamp 1676037725
transform 1 0 4232 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_46
timestamp 1676037725
transform 1 0 5336 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_8
timestamp 1676037725
transform 1 0 1840 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_33
timestamp 1676037725
transform 1 0 4140 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_40
timestamp 1676037725
transform 1 0 4784 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_9
timestamp 1676037725
transform 1 0 1932 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_17
timestamp 1676037725
transform 1 0 2668 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_21
timestamp 1676037725
transform 1 0 3036 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1676037725
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_34
timestamp 1676037725
transform 1 0 4232 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_47
timestamp 1676037725
transform 1 0 5428 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_9
timestamp 1676037725
transform 1 0 1932 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_19
timestamp 1676037725
transform 1 0 2852 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_40
timestamp 1676037725
transform 1 0 4784 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_7
timestamp 1676037725
transform 1 0 1748 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_11
timestamp 1676037725
transform 1 0 2116 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1676037725
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_45
timestamp 1676037725
transform 1 0 5244 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_7
timestamp 1676037725
transform 1 0 1748 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_11
timestamp 1676037725
transform 1 0 2116 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_36
timestamp 1676037725
transform 1 0 4416 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_46
timestamp 1676037725
transform 1 0 5336 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_11
timestamp 1676037725
transform 1 0 2116 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_20
timestamp 1676037725
transform 1 0 2944 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_37
timestamp 1676037725
transform 1 0 4508 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_43
timestamp 1676037725
transform 1 0 5060 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_47
timestamp 1676037725
transform 1 0 5428 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_23
timestamp 1676037725
transform 1 0 3220 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_46
timestamp 1676037725
transform 1 0 5336 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_47
timestamp 1676037725
transform 1 0 5428 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_9
timestamp 1676037725
transform 1 0 1932 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_21
timestamp 1676037725
transform 1 0 3036 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_33
timestamp 1676037725
transform 1 0 4140 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_41
timestamp 1676037725
transform 1 0 4876 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_46
timestamp 1676037725
transform 1 0 5336 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_9
timestamp 1676037725
transform 1 0 1932 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_20
timestamp 1676037725
transform 1 0 2944 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_35
timestamp 1676037725
transform 1 0 4324 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_46
timestamp 1676037725
transform 1 0 5336 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 5796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 5796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 5796 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 5796 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 5796 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 5796 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 5796 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 5796 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 5796 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 5796 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 5796 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 5796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 5796 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__and3_1  _11_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2484 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _12_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2300 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _13_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4600 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _14_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3956 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _15_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2116 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _16_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 2116 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _17_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2024 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _18_
timestamp 1676037725
transform -1 0 5244 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _19_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2852 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _20_
timestamp 1676037725
transform 1 0 3956 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _21_
timestamp 1676037725
transform -1 0 1840 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _22_
timestamp 1676037725
transform -1 0 5060 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _23_
timestamp 1676037725
transform -1 0 4784 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _24_
timestamp 1676037725
transform -1 0 4232 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _25_
timestamp 1676037725
transform -1 0 4876 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _26_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3496 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _27_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2208 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _28_
timestamp 1676037725
transform 1 0 3496 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _29_
timestamp 1676037725
transform -1 0 3496 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2944 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1676037725
transform -1 0 3496 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1676037725
transform 1 0 2576 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2024 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform -1 0 5336 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4968 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp 1676037725
transform -1 0 2668 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 1676037725
transform 1 0 4968 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1676037725
transform -1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1676037725
transform -1 0 1932 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1676037725
transform 1 0 4968 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1676037725
transform 1 0 3128 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1676037725
transform -1 0 1932 0 -1 8704
box -38 -48 406 592
<< labels >>
flabel metal4 s 2604 2128 2924 9296 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 1944 2128 2264 9296 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 clk
port 2 nsew signal input
flabel metal3 s 6100 2728 6900 2848 0 FreeSans 480 0 0 0 counter[0]
port 3 nsew signal tristate
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 counter[1]
port 4 nsew signal tristate
flabel metal2 s 5170 10624 5226 11424 0 FreeSans 224 90 0 0 counter[2]
port 5 nsew signal tristate
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 counter[3]
port 6 nsew signal tristate
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 countern[0]
port 7 nsew signal tristate
flabel metal3 s 6100 9528 6900 9648 0 FreeSans 480 0 0 0 countern[1]
port 8 nsew signal tristate
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 countern[2]
port 9 nsew signal tristate
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 countern[3]
port 10 nsew signal tristate
flabel metal2 s 1950 10624 2006 11424 0 FreeSans 224 90 0 0 en
port 11 nsew signal input
flabel metal3 s 6100 6128 6900 6248 0 FreeSans 480 0 0 0 reset
port 12 nsew signal input
rlabel metal1 3450 8704 3450 8704 0 VGND
rlabel metal1 3450 9248 3450 9248 0 VPWR
rlabel metal2 4922 7106 4922 7106 0 _00_
rlabel metal1 4646 4148 4646 4148 0 _01_
rlabel metal2 4278 3230 4278 3230 0 _02_
rlabel metal1 2070 3543 2070 3543 0 _03_
rlabel metal1 3634 5814 3634 5814 0 _04_
rlabel metal1 2576 2958 2576 2958 0 _05_
rlabel metal2 3818 4318 3818 4318 0 _06_
rlabel metal1 3910 3434 3910 3434 0 _07_
rlabel metal1 2300 5066 2300 5066 0 _08_
rlabel metal1 4002 5746 4002 5746 0 _09_
rlabel metal2 2944 6324 2944 6324 0 _10_
rlabel metal3 820 6868 820 6868 0 clk
rlabel metal1 4186 5338 4186 5338 0 clknet_0_clk
rlabel metal2 3542 2788 3542 2788 0 clknet_1_0__leaf_clk
rlabel metal2 3910 4998 3910 4998 0 clknet_1_1__leaf_clk
rlabel metal1 5336 2618 5336 2618 0 counter[0]
rlabel metal2 46 2744 46 2744 0 counter[1]
rlabel metal2 5198 9904 5198 9904 0 counter[2]
rlabel metal2 6486 1520 6486 1520 0 counter[3]
rlabel metal3 820 3468 820 3468 0 countern[0]
rlabel metal1 5566 8602 5566 8602 0 countern[1]
rlabel metal2 3266 2608 3266 2608 0 countern[2]
rlabel metal1 1334 8602 1334 8602 0 countern[3]
rlabel metal1 1978 9010 1978 9010 0 en
rlabel metal2 2438 4148 2438 4148 0 net1
rlabel metal1 3082 5712 3082 5712 0 net10
rlabel metal2 4738 3808 4738 3808 0 net2
rlabel metal1 4508 3910 4508 3910 0 net3
rlabel metal2 4002 3876 4002 3876 0 net4
rlabel metal1 3358 6834 3358 6834 0 net5
rlabel metal1 4876 5678 4876 5678 0 net6
rlabel metal2 1886 5338 1886 5338 0 net7
rlabel metal1 4554 4794 4554 4794 0 net8
rlabel metal1 1932 4046 1932 4046 0 net9
rlabel metal1 5566 6290 5566 6290 0 reset
<< properties >>
string FIXED_BBOX 0 0 6900 11424
<< end >>
