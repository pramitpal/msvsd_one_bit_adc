magic
tech sky130A
magscale 1 2
timestamp 1678560175
<< error_p >>
rect 2183 2732 2202 2752
<< metal3 >>
rect 53 2732 2183 2852
rect 53 2692 2232 2732
rect 2142 2534 2232 2692
rect 172 474 2232 2534
rect 53 284 2183 332
rect 53 220 230 284
rect 294 220 2183 284
rect 53 172 2183 220
<< via3 >>
rect 230 220 294 284
<< mimcap >>
rect 202 616 2202 2504
rect 202 552 230 616
rect 294 552 2202 616
rect 202 504 2202 552
<< mimcapcontact >>
rect 230 552 294 616
<< metal4 >>
rect 217 616 307 670
rect 217 552 230 616
rect 294 552 307 616
rect 217 284 307 552
rect 217 220 230 284
rect 294 220 307 284
rect 217 166 307 220
<< end >>
