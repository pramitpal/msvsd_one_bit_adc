magic
tech sky130A
magscale 1 2
timestamp 1677774298
<< nwell >>
rect 188 178 616 386
<< nmos >>
rect 282 -12 312 72
rect 492 -12 522 72
<< pmos >>
rect 282 240 312 324
rect 492 240 522 324
<< ndiff >>
rect 224 60 282 72
rect 224 0 236 60
rect 270 0 282 60
rect 224 -12 282 0
rect 312 60 370 72
rect 312 0 324 60
rect 358 0 370 60
rect 312 -12 370 0
rect 434 60 492 72
rect 434 0 446 60
rect 480 0 492 60
rect 434 -12 492 0
rect 522 60 580 72
rect 522 0 534 60
rect 568 0 580 60
rect 522 -12 580 0
<< pdiff >>
rect 224 312 282 324
rect 224 252 236 312
rect 270 252 282 312
rect 224 240 282 252
rect 312 312 370 324
rect 312 252 324 312
rect 358 252 370 312
rect 312 240 370 252
rect 434 312 492 324
rect 434 252 446 312
rect 480 252 492 312
rect 434 240 492 252
rect 522 312 580 324
rect 522 252 534 312
rect 568 252 580 312
rect 522 240 580 252
<< ndiffc >>
rect 236 0 270 60
rect 324 0 358 60
rect 446 0 480 60
rect 534 0 568 60
<< pdiffc >>
rect 236 252 270 312
rect 324 252 358 312
rect 446 252 480 312
rect 534 252 568 312
<< poly >>
rect 282 324 312 350
rect 492 324 522 350
rect -27 159 27 175
rect -27 125 -17 159
rect 17 157 27 159
rect 70 157 100 237
rect 17 127 100 157
rect 17 125 27 127
rect -27 109 27 125
rect 70 80 100 127
rect 173 159 239 169
rect 173 125 189 159
rect 223 157 239 159
rect 282 157 312 240
rect 223 127 312 157
rect 223 125 239 127
rect 173 115 239 125
rect 282 72 312 127
rect 383 159 449 169
rect 383 125 399 159
rect 433 157 449 159
rect 492 157 522 240
rect 433 127 522 157
rect 433 125 449 127
rect 383 115 449 125
rect 492 72 522 127
rect 282 -38 312 -12
rect 492 -38 522 -12
<< polycont >>
rect -17 125 17 159
rect 189 125 223 159
rect 399 125 433 159
<< locali >>
rect 236 312 270 328
rect 236 236 270 252
rect 324 312 358 328
rect 324 236 358 252
rect 446 312 480 328
rect 446 236 480 252
rect 534 312 568 328
rect 534 236 568 252
rect 189 159 223 175
rect -33 125 -17 159
rect 17 125 33 159
rect 189 109 223 125
rect 399 159 433 175
rect 399 109 433 125
rect 236 60 270 76
rect 236 -16 270 0
rect 324 60 358 76
rect 324 -16 358 0
rect 446 60 480 76
rect 446 -16 480 0
rect 534 60 568 76
rect 534 -16 568 0
<< viali >>
rect 236 252 270 312
rect 324 252 358 312
rect 446 252 480 312
rect 534 252 568 312
rect -17 125 17 159
rect 189 125 223 159
rect 399 125 433 159
rect 236 0 270 60
rect 324 0 358 60
rect 446 0 480 60
rect 534 0 568 60
<< metal1 >>
rect 24 435 58 437
rect 24 431 267 435
rect 24 401 479 431
rect 24 310 58 401
rect 233 397 479 401
rect 233 324 267 397
rect 445 324 479 397
rect 230 312 276 324
rect 230 252 236 312
rect 270 252 276 312
rect -26 168 26 174
rect -29 119 -26 165
rect 26 119 29 165
rect 114 159 146 252
rect 230 240 276 252
rect 318 312 364 324
rect 318 252 324 312
rect 358 252 364 312
rect 318 240 364 252
rect 440 312 486 324
rect 440 252 446 312
rect 480 252 486 312
rect 440 240 486 252
rect 528 312 574 324
rect 528 252 534 312
rect 568 252 574 312
rect 528 240 574 252
rect 183 159 229 171
rect 114 125 189 159
rect 223 125 229 159
rect -26 110 26 116
rect 114 66 146 125
rect 183 113 229 125
rect 326 159 358 240
rect 393 159 439 171
rect 326 125 399 159
rect 433 125 439 159
rect 326 72 358 125
rect 393 113 439 125
rect 536 159 568 240
rect 596 168 648 174
rect 536 125 596 159
rect 536 72 568 125
rect 596 110 648 116
rect 230 60 276 72
rect 26 -69 60 18
rect 230 0 236 60
rect 270 0 276 60
rect 230 -12 276 0
rect 318 60 364 72
rect 318 0 324 60
rect 358 0 364 60
rect 318 -12 364 0
rect 440 60 486 72
rect 440 0 446 60
rect 480 0 486 60
rect 440 -12 486 0
rect 528 60 574 72
rect 528 0 534 60
rect 568 0 574 60
rect 528 -12 574 0
rect 237 -65 271 -12
rect 451 -65 485 -12
rect 237 -69 485 -65
rect 26 -99 485 -69
rect 26 -103 271 -99
<< via1 >>
rect -26 159 26 168
rect -26 125 -17 159
rect -17 125 17 159
rect 17 125 26 159
rect -26 116 26 125
rect 596 116 648 168
<< metal2 >>
rect -32 116 -26 168
rect 26 159 32 168
rect 590 159 596 168
rect 26 125 596 159
rect 26 116 32 125
rect 590 116 596 125
rect 648 116 654 168
use sky130_fd_pr__nfet_01v8_KMMFGM  sky130_fd_pr__nfet_01v8_KMMFGM_0
timestamp 1677774298
transform 1 0 85 0 1 30
box -73 -68 73 68
use sky130_fd_pr__pfet_01v8_2ZVT9K  sky130_fd_pr__pfet_01v8_2ZVT9K_0
timestamp 1677774298
transform 1 0 85 0 1 282
box -109 -104 109 104
<< labels >>
flabel metal1 s 252 412 252 412 3 FreeSans 800 0 0 0 VDD
flabel metal2 s 620 140 620 140 3 FreeSans 800 0 0 0 Y
flabel metal1 s 256 -78 256 -78 3 FreeSans 800 0 0 0 GND
<< end >>
