* SPICE3 file created from RING_OSC_0.ext - technology: sky130A

X0 m1_688_4424# li_405_1579# m1_398_2912# m1_398_2912# sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.12 as=0.2226 ps=2.21 w=0.84 l=0.15
X1 m1_398_2912# li_405_1579# m1_688_4424# m1_398_2912# sky130_fd_pr__pfet_01v8 ad=0.2226 pd=2.21 as=0.1176 ps=1.12 w=0.84 l=0.15
X2 m1_688_4424# li_405_1579# SUB SUB sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2226 ps=2.21 w=0.84 l=0.15
X3 SUB li_405_1579# m1_688_4424# SUB sky130_fd_pr__nfet_01v8 ad=0.2226 pd=2.21 as=0.1176 ps=1.12 w=0.84 l=0.15
X4 STAGE2_INV_48448484_0_0_1677766866_0/li_491_571# m1_688_4424# m1_398_2912# m1_398_2912# sky130_fd_pr__pfet_01v8 ad=0.1176 pd=1.12 as=0.2226 ps=2.21 w=0.84 l=0.15
X5 m1_398_2912# m1_688_4424# STAGE2_INV_48448484_0_0_1677766866_0/li_491_571# m1_398_2912# sky130_fd_pr__pfet_01v8 ad=0.2226 pd=2.21 as=0.1176 ps=1.12 w=0.84 l=0.15
X6 li_405_1579# STAGE2_INV_48448484_0_0_1677766866_0/li_491_571# m1_398_2912# m1_398_2912# sky130_fd_pr__pfet_01v8 ad=0.2352 pd=2.24 as=1.3356 ps=13.26 w=0.84 l=0.15
X7 m1_398_2912# STAGE2_INV_48448484_0_0_1677766866_0/li_491_571# li_405_1579# m1_398_2912# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
X8 li_405_1579# STAGE2_INV_48448484_0_0_1677766866_0/li_491_571# SUB SUB sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2226 ps=2.21 w=0.84 l=0.15
X9 SUB STAGE2_INV_48448484_0_0_1677766866_0/li_491_571# li_405_1579# SUB sky130_fd_pr__nfet_01v8 ad=0.2226 pd=2.21 as=0.1176 ps=1.12 w=0.84 l=0.15
X10 STAGE2_INV_48448484_0_0_1677766866_0/li_491_571# m1_688_4424# SUB SUB sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.24 as=1.3356 ps=13.26 w=0.84 l=0.15
X11 SUB m1_688_4424# STAGE2_INV_48448484_0_0_1677766866_0/li_491_571# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.84 l=0.15
