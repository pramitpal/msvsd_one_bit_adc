magic
tech sky130A
magscale 1 2
timestamp 1678560175
<< locali >>
rect 1695 6955 1703 6989
rect 1737 6955 1745 6989
rect 1695 6905 1745 6955
rect 1695 6871 1703 6905
rect 1737 6871 1745 6905
rect 577 6031 585 6065
rect 619 6031 627 6065
rect 577 5981 627 6031
rect 577 5947 585 5981
rect 619 5947 627 5981
rect 1437 5107 1445 5141
rect 1479 5107 1487 5141
rect 1437 5057 1487 5107
rect 1437 5023 1445 5057
rect 1479 5023 1487 5057
rect 2813 4435 2821 4469
rect 2855 4435 2863 4469
rect 2813 3965 2863 4435
rect 2813 3931 2821 3965
rect 2855 3931 2863 3965
<< viali >>
rect 1703 6955 1737 6989
rect 1703 6871 1737 6905
rect 585 6031 619 6065
rect 585 5947 619 5981
rect 1445 5107 1479 5141
rect 1445 5023 1479 5057
rect 2821 4435 2855 4469
rect 2821 3931 2855 3965
<< metal1 >>
rect 1686 6989 1978 7000
rect 1686 6955 1703 6989
rect 1737 6955 1978 6989
rect 1686 6944 1978 6955
rect 1258 6914 1754 6916
rect 1258 6862 1264 6914
rect 1316 6905 1754 6914
rect 1316 6871 1703 6905
rect 1737 6871 1754 6905
rect 1316 6862 1754 6871
rect 1258 6860 1754 6862
rect 2032 6326 2182 6328
rect 2032 6274 2038 6326
rect 2090 6274 2124 6326
rect 2176 6274 2182 6326
rect 2032 6272 2182 6274
rect 1000 6242 1118 6244
rect 1000 6190 1006 6242
rect 1058 6190 1118 6242
rect 1000 6188 1118 6190
rect 1860 6158 1978 6160
rect 1860 6106 1866 6158
rect 1918 6106 1978 6158
rect 1860 6104 1978 6106
rect 226 6074 636 6076
rect 226 6022 232 6074
rect 284 6065 636 6074
rect 284 6031 585 6065
rect 619 6031 636 6065
rect 284 6022 636 6031
rect 226 6020 636 6022
rect 357 5936 478 5992
rect 568 5981 946 5992
rect 568 5947 585 5981
rect 619 5947 946 5981
rect 568 5936 946 5947
rect 1000 5990 1064 5992
rect 1000 5938 1006 5990
rect 1058 5938 1064 5990
rect 1000 5936 1064 5938
rect 1258 5990 1634 5992
rect 1258 5938 1264 5990
rect 1316 5938 1634 5990
rect 1258 5936 1634 5938
rect 1172 5906 1236 5908
rect 1172 5854 1178 5906
rect 1230 5854 1236 5906
rect 1172 5852 1236 5854
rect 1516 5906 1580 5908
rect 1516 5854 1522 5906
rect 1574 5854 1580 5906
rect 1516 5852 1580 5854
rect 1860 5906 1924 5908
rect 1860 5854 1866 5906
rect 1918 5854 1924 5906
rect 1860 5852 1924 5854
rect 1172 5822 1580 5824
rect 1172 5770 1178 5822
rect 1230 5770 1522 5822
rect 1574 5770 1580 5822
rect 1172 5768 1580 5770
rect 2634 5318 3214 5320
rect 2634 5266 2640 5318
rect 2692 5266 3156 5318
rect 3208 5266 3214 5318
rect 2634 5264 3214 5266
rect 1118 5141 1496 5152
rect 1118 5107 1445 5141
rect 1479 5107 1496 5141
rect 1118 5096 1496 5107
rect 1694 5096 1750 5184
rect 1428 5066 2354 5068
rect 1428 5057 2296 5066
rect 1428 5023 1445 5057
rect 1479 5023 2296 5057
rect 1428 5014 2296 5023
rect 2348 5014 2354 5066
rect 1428 5012 2354 5014
rect 2462 4814 2784 4816
rect 2462 4762 2468 4814
rect 2520 4762 2726 4814
rect 2778 4762 2784 4814
rect 2462 4760 2784 4762
rect 914 4730 978 4732
rect 914 4678 920 4730
rect 972 4678 978 4730
rect 914 4676 978 4678
rect 1602 4730 1666 4732
rect 1602 4678 1608 4730
rect 1660 4678 1666 4730
rect 1602 4676 1666 4678
rect 2494 4478 2698 4480
rect 2494 4426 2640 4478
rect 2692 4426 2698 4478
rect 2494 4424 2698 4426
rect 2804 4478 3010 4480
rect 2804 4426 2812 4478
rect 2864 4426 3010 4478
rect 2804 4424 3010 4426
rect 3182 4424 3698 4480
rect 2204 4310 2526 4312
rect 2204 4258 2210 4310
rect 2262 4258 2468 4310
rect 2520 4258 2526 4310
rect 2204 4256 2526 4258
rect 1118 3920 1634 3976
rect 1806 3965 2872 3976
rect 1806 3931 2821 3965
rect 2855 3931 2872 3965
rect 1806 3920 2872 3931
rect 2204 3638 2322 3640
rect 2204 3586 2210 3638
rect 2262 3586 2322 3638
rect 2204 3584 2322 3586
rect 2634 3638 3042 3640
rect 2634 3586 2640 3638
rect 2692 3586 2984 3638
rect 3036 3586 3042 3638
rect 2634 3584 3042 3586
rect 3182 3584 3698 3640
rect 1000 3134 1064 3136
rect 1000 3082 1006 3134
rect 1058 3082 1064 3134
rect 1000 3080 1064 3082
rect 1602 3134 1666 3136
rect 1602 3082 1608 3134
rect 1660 3082 1666 3134
rect 1602 3080 1666 3082
<< via1 >>
rect 1264 6862 1316 6914
rect 2038 6274 2090 6326
rect 2124 6274 2176 6326
rect 1006 6190 1058 6242
rect 1866 6106 1918 6158
rect 232 6022 284 6074
rect 1006 5938 1058 5990
rect 1264 5938 1316 5990
rect 1178 5854 1230 5906
rect 1522 5854 1574 5906
rect 1866 5854 1918 5906
rect 1178 5770 1230 5822
rect 1522 5770 1574 5822
rect 2640 5266 2692 5318
rect 3156 5266 3208 5318
rect 2296 5014 2348 5066
rect 2468 4762 2520 4814
rect 2726 4762 2778 4814
rect 920 4678 972 4730
rect 1608 4678 1660 4730
rect 2640 4426 2692 4478
rect 2812 4469 2864 4478
rect 2812 4435 2821 4469
rect 2821 4435 2855 4469
rect 2855 4435 2864 4469
rect 2812 4426 2864 4435
rect 2210 4258 2262 4310
rect 2468 4258 2520 4310
rect 2210 3586 2262 3638
rect 2640 3586 2692 3638
rect 2984 3586 3036 3638
rect 1006 3082 1058 3134
rect 1608 3082 1660 3134
<< metal2 >>
rect 2724 7336 2780 7345
rect 402 7084 458 7093
rect 402 7019 458 7028
rect 1090 7084 1146 7093
rect 1090 7019 1146 7028
rect 1262 6914 1318 6920
rect 1262 6862 1264 6914
rect 1316 6862 1318 6914
rect 1262 6856 1318 6862
rect 2036 6326 2092 6332
rect 2036 6274 2038 6326
rect 2090 6274 2092 6326
rect 1004 6242 1060 6248
rect 1004 6190 1006 6242
rect 1058 6190 1060 6242
rect 230 6074 286 6080
rect 230 6022 232 6074
rect 284 6022 286 6074
rect 230 6016 286 6022
rect 1004 5990 1060 6190
rect 1864 6158 1920 6164
rect 1004 5938 1006 5990
rect 1058 5938 1060 5990
rect 1004 5932 1060 5938
rect 1262 5990 1318 6132
rect 1262 5938 1264 5990
rect 1316 5938 1318 5990
rect 1262 5932 1318 5938
rect 1864 6106 1866 6158
rect 1918 6106 1920 6158
rect 1176 5906 1232 5912
rect 1176 5854 1178 5906
rect 1230 5854 1232 5906
rect 1176 5822 1232 5854
rect 1176 5770 1178 5822
rect 1230 5770 1232 5822
rect 1176 5764 1232 5770
rect 1520 5906 1576 5912
rect 1520 5854 1522 5906
rect 1574 5854 1576 5906
rect 1520 5822 1576 5854
rect 1864 5906 1920 6106
rect 1864 5854 1866 5906
rect 1918 5854 1920 5906
rect 1864 5848 1920 5854
rect 1520 5770 1522 5822
rect 1574 5770 1576 5822
rect 1520 5764 1576 5770
rect 144 5320 200 5329
rect 144 280 200 5264
rect 402 5320 458 5329
rect 402 5255 458 5264
rect 918 5320 974 5329
rect 918 4730 974 5264
rect 918 4678 920 4730
rect 972 4678 974 4730
rect 918 4672 974 4678
rect 1606 5320 1662 5329
rect 1606 4730 1662 5264
rect 1606 4678 1608 4730
rect 1660 4678 1662 4730
rect 1606 4672 1662 4678
rect 1778 5320 1834 5329
rect 1778 4368 1834 5264
rect 2036 5320 2092 6274
rect 2122 6326 2178 6332
rect 2122 6274 2124 6326
rect 2176 6274 2178 6326
rect 2122 6268 2178 6274
rect 2036 5255 2092 5264
rect 2208 5320 2264 5329
rect 2208 4310 2264 5264
rect 2552 5320 2608 5329
rect 2294 5066 2350 5072
rect 2294 5014 2296 5066
rect 2348 5014 2350 5066
rect 2294 5008 2350 5014
rect 2466 4814 2522 4820
rect 2466 4762 2468 4814
rect 2520 4762 2522 4814
rect 2466 4756 2522 4762
rect 2208 4258 2210 4310
rect 2262 4258 2264 4310
rect 2208 4252 2264 4258
rect 2466 4310 2522 4316
rect 2466 4258 2468 4310
rect 2520 4258 2522 4310
rect 2466 4252 2522 4258
rect 2208 3638 2264 3644
rect 2208 3586 2210 3638
rect 2262 3586 2264 3638
rect 1090 3556 1146 3565
rect 1090 3491 1146 3500
rect 1004 3134 1060 3140
rect 1004 3082 1006 3134
rect 1058 3082 1060 3134
rect 1004 2800 1060 3082
rect 1004 2735 1060 2744
rect 1606 3134 1662 3140
rect 1606 3082 1608 3134
rect 1660 3082 1662 3134
rect 1606 2800 1662 3082
rect 1606 2735 1662 2744
rect 2208 2800 2264 3586
rect 2208 2735 2264 2744
rect 144 215 200 224
rect 2552 280 2608 5264
rect 2638 5320 2694 5329
rect 2638 5255 2694 5264
rect 2724 5320 2780 7280
rect 2724 5255 2780 5264
rect 3154 5318 3210 5324
rect 3154 5266 3156 5318
rect 3208 5266 3210 5318
rect 2724 4814 2780 4820
rect 2724 4762 2726 4814
rect 2778 4762 2780 4814
rect 2638 4478 2694 4484
rect 2638 4426 2640 4478
rect 2692 4426 2694 4478
rect 2638 3638 2694 4426
rect 2638 3586 2640 3638
rect 2692 3586 2694 3638
rect 2638 3580 2694 3586
rect 2724 3556 2780 4762
rect 2810 4816 2866 4825
rect 2810 4478 2866 4760
rect 2810 4426 2812 4478
rect 2864 4426 2866 4478
rect 2810 4420 2866 4426
rect 3154 4368 3210 5266
rect 2724 3491 2780 3500
rect 2982 3638 3038 3644
rect 2982 3586 2984 3638
rect 3036 3586 3038 3638
rect 2982 2800 3038 3586
rect 3842 3556 3898 3565
rect 3842 3491 3898 3500
rect 2982 2735 3038 2744
rect 2552 215 2608 224
<< via2 >>
rect 2724 7280 2780 7336
rect 402 7028 458 7084
rect 1090 7028 1146 7084
rect 144 5264 200 5320
rect 402 5264 458 5320
rect 918 5264 974 5320
rect 1606 5264 1662 5320
rect 1778 5264 1834 5320
rect 2036 5264 2092 5320
rect 2208 5264 2264 5320
rect 2552 5264 2608 5320
rect 1090 3500 1146 3556
rect 1004 2744 1060 2800
rect 1606 2744 1662 2800
rect 2208 2744 2264 2800
rect 144 224 200 280
rect 2638 5318 2694 5320
rect 2638 5266 2640 5318
rect 2640 5266 2692 5318
rect 2692 5266 2694 5318
rect 2638 5264 2694 5266
rect 2724 5264 2780 5320
rect 2810 4760 2866 4816
rect 2724 3500 2780 3556
rect 3842 3500 3898 3556
rect 2982 2744 3038 2800
rect 2552 224 2608 280
<< metal3 >>
rect 2719 7336 2838 7388
rect 2719 7280 2724 7336
rect 2780 7280 2838 7336
rect 2719 7228 2838 7280
rect -80 7088 2832 7136
rect -80 7084 2336 7088
rect -80 7028 402 7084
rect 458 7028 1090 7084
rect 1146 7028 2336 7084
rect -80 7024 2336 7028
rect 2400 7024 2832 7088
rect -80 6976 2832 7024
rect -80 5324 2832 5372
rect -80 5260 -32 5324
rect 32 5320 2832 5324
rect 32 5264 144 5320
rect 200 5264 402 5320
rect 458 5264 918 5320
rect 974 5264 1606 5320
rect 1662 5264 1778 5320
rect 1834 5264 2036 5320
rect 2092 5264 2208 5320
rect 2264 5264 2552 5320
rect 2608 5264 2638 5320
rect 2694 5264 2724 5320
rect 2780 5264 2832 5320
rect 32 5260 2832 5264
rect -80 5212 2832 5260
rect 2805 4816 2871 4868
rect 2805 4760 2810 4816
rect 2866 4760 2871 4816
rect 2805 4708 2871 4760
rect 4894 4713 4984 4983
rect -80 3560 4896 3608
rect -80 3556 2336 3560
rect -80 3500 1090 3556
rect 1146 3500 2336 3556
rect -80 3496 2336 3500
rect 2400 3556 4896 3560
rect 2400 3500 2724 3556
rect 2780 3500 3842 3556
rect 3898 3500 4896 3556
rect 2400 3496 4896 3500
rect -80 3448 4896 3496
rect 90 2581 180 2851
rect 999 2800 1065 2852
rect 999 2744 1004 2800
rect 1060 2744 1065 2800
rect 999 2692 1065 2744
rect 1601 2800 1667 2852
rect 1601 2744 1606 2800
rect 1662 2744 1667 2800
rect 1601 2692 1667 2744
rect 2203 2800 2269 2852
rect 2203 2744 2208 2800
rect 2264 2744 2269 2800
rect 2203 2692 2269 2744
rect 2977 2800 3043 2852
rect 2977 2744 2982 2800
rect 3038 2744 3043 2800
rect 2977 2692 3043 2744
rect 4464 2589 4554 2841
rect 139 280 205 332
rect 139 224 144 280
rect 200 224 205 280
rect 139 172 205 224
rect 2547 280 2613 332
rect 2547 224 2552 280
rect 2608 224 2613 280
rect 2547 172 2613 224
<< via3 >>
rect 2336 7024 2400 7088
rect -32 5260 32 5324
rect 2336 3496 2400 3560
<< metal4 >>
rect -118 5324 118 7174
rect -118 5260 -32 5324
rect 32 5260 118 5324
rect -118 -118 118 5260
rect 2250 7088 2486 7174
rect 2250 7024 2336 7088
rect 2400 7024 2486 7088
rect 2250 3560 2486 7024
rect 2250 3496 2336 3560
rect 2400 3496 2486 3560
rect 2250 1646 2486 3496
use CAP_2T_51284459_1678559787  CAP_2T_51284459_1678559787_0
timestamp 1678560175
transform -1 0 2322 0 1 0
box 53 166 2232 2852
use CAP_2T_51284459_1678559787  CAP_2T_51284459_1678559787_1
timestamp 1678560175
transform 1 0 2752 0 -1 7560
box 53 166 2232 2852
use CAP_2T_51284459_1678559787  CAP_2T_51284459_1678559787_2
timestamp 1678560175
transform 1 0 2322 0 1 0
box 53 166 2232 2852
use INV_97143719_PG0_0_0_1678559785  INV_97143719_PG0_0_0_1678559785_0
timestamp 1678560175
transform 1 0 0 0 1 4536
box 0 30 688 3024
use INV_97143719_PG0_1_0_1678559786  INV_97143719_PG0_1_0_1678559786_0
timestamp 1678560175
transform 1 0 2064 0 1 3024
box 0 30 688 3024
use NMOS_4T_41917219_X2_Y1_1678559788  NMOS_4T_41917219_X2_Y1_1678559788_0
timestamp 1678560175
transform 1 0 1376 0 -1 6048
box 121 56 567 1482
use NMOS_4T_41917219_X2_Y1_1678559788  NMOS_4T_41917219_X2_Y1_1678559788_1
timestamp 1678560175
transform 1 0 688 0 -1 6048
box 121 56 567 1482
use NMOS_S_97312901_X2_Y1_1678559789  NMOS_S_97312901_X2_Y1_1678559789_0
timestamp 1678560175
transform 1 0 1720 0 1 6048
box 121 56 567 1482
use NMOS_S_97312901_X2_Y1_1678559789  NMOS_S_97312901_X2_Y1_1678559789_1
timestamp 1678560175
transform 1 0 1376 0 1 3024
box 121 56 567 1482
use NMOS_S_97312901_X2_Y1_1678559789  NMOS_S_97312901_X2_Y1_1678559789_2
timestamp 1678560175
transform 1 0 2752 0 -1 4536
box 121 56 567 1482
use PMOS_S_78930897_X2_Y1_1678559790  PMOS_S_78930897_X2_Y1_1678559790_0
timestamp 1678560175
transform 1 0 688 0 1 3024
box 0 0 688 1512
use PMOS_S_78930897_X2_Y1_1678559790  PMOS_S_78930897_X2_Y1_1678559790_1
timestamp 1678560175
transform 1 0 3440 0 -1 4536
box 0 0 688 1512
use SCM_PMOS_79287875_X2_Y1_1678559791  SCM_PMOS_79287875_X2_Y1_1678559791_0
timestamp 1678560175
transform -1 0 1720 0 1 6048
box 0 0 1032 1512
<< labels >>
flabel metal3 s 1204 2772 1204 2772 0 FreeSerif 0 0 0 0 INP
port 2 nsew
flabel metal4 s 0 4410 0 4410 0 FreeSerif 0 0 0 0 GND
port 4 nsew
flabel metal2 s 2580 2772 2580 2772 0 FreeSerif 0 0 0 0 GND
port 4 nsew
flabel metal4 s 0 4410 0 4410 0 FreeSerif 0 0 0 0 GND
port 4 nsew
flabel metal4 s 0 4410 0 4410 0 FreeSerif 0 0 0 0 GND
port 4 nsew
flabel metal4 s 0 4410 0 4410 0 FreeSerif 0 0 0 0 GND
port 4 nsew
flabel metal4 s 0 4410 0 4410 0 FreeSerif 0 0 0 0 GND
port 4 nsew
flabel metal4 s 0 4410 0 4410 0 FreeSerif 0 0 0 0 GND
port 4 nsew
flabel metal4 s 0 4410 0 4410 0 FreeSerif 0 0 0 0 GND
port 4 nsew
flabel metal4 s 0 4410 0 4410 0 FreeSerif 0 0 0 0 GND
port 4 nsew
flabel metal4 s 0 4410 0 4410 0 FreeSerif 0 0 0 0 GND
port 4 nsew
flabel metal4 s 0 4410 0 4410 0 FreeSerif 0 0 0 0 GND
port 4 nsew
flabel metal4 s 0 4410 0 4410 0 FreeSerif 0 0 0 0 GND
port 4 nsew
flabel metal4 s 0 4410 0 4410 0 FreeSerif 0 0 0 0 GND
port 4 nsew
flabel metal4 s 0 4410 0 4410 0 FreeSerif 0 0 0 0 GND
port 4 nsew
flabel metal4 s 0 4410 0 4410 0 FreeSerif 0 0 0 0 GND
port 4 nsew
flabel metal4 s 0 4410 0 4410 0 FreeSerif 0 0 0 0 GND
port 4 nsew
flabel metal4 s 0 4410 0 4410 0 FreeSerif 0 0 0 0 GND
port 4 nsew
flabel metal4 s 0 4410 0 4410 0 FreeSerif 0 0 0 0 GND
port 4 nsew
flabel metal4 s 0 4410 0 4410 0 FreeSerif 0 0 0 0 GND
port 4 nsew
flabel metal4 s 0 4410 0 4410 0 FreeSerif 0 0 0 0 GND
port 4 nsew
flabel metal4 s 0 4410 0 4410 0 FreeSerif 0 0 0 0 GND
port 4 nsew
flabel metal4 s 0 4410 0 4410 0 FreeSerif 0 0 0 0 GND
port 4 nsew
flabel metal4 s 0 4410 0 4410 0 FreeSerif 0 0 0 0 GND
port 4 nsew
flabel metal4 s 0 4410 0 4410 0 FreeSerif 0 0 0 0 GND
port 4 nsew
flabel metal4 s 0 4410 0 4410 0 FreeSerif 0 0 0 0 GND
port 4 nsew
flabel metal4 s 0 4410 0 4410 0 FreeSerif 0 0 0 0 GND
port 4 nsew
flabel metal4 s 0 4410 0 4410 0 FreeSerif 0 0 0 0 GND
port 4 nsew
flabel metal4 s 0 4410 0 4410 0 FreeSerif 0 0 0 0 GND
port 4 nsew
flabel metal4 s 0 4410 0 4410 0 FreeSerif 0 0 0 0 GND
port 4 nsew
flabel metal4 s 0 4410 0 4410 0 FreeSerif 0 0 0 0 GND
port 4 nsew
flabel metal4 s 0 4410 0 4410 0 FreeSerif 0 0 0 0 GND
port 4 nsew
flabel metal4 s 0 4410 0 4410 0 FreeSerif 0 0 0 0 GND
port 4 nsew
flabel metal4 s 2368 4410 2368 4410 0 FreeSerif 0 0 0 0 VDD
port 5 nsew
flabel metal4 s 2368 4410 2368 4410 0 FreeSerif 0 0 0 0 VDD
port 5 nsew
flabel metal4 s 2368 4410 2368 4410 0 FreeSerif 0 0 0 0 VDD
port 5 nsew
flabel metal4 s 2368 4410 2368 4410 0 FreeSerif 0 0 0 0 VDD
port 5 nsew
flabel metal4 s 2368 4410 2368 4410 0 FreeSerif 0 0 0 0 VDD
port 5 nsew
flabel metal4 s 2368 4410 2368 4410 0 FreeSerif 0 0 0 0 VDD
port 5 nsew
flabel metal4 s 2368 4410 2368 4410 0 FreeSerif 0 0 0 0 VDD
port 5 nsew
flabel metal4 s 2368 4410 2368 4410 0 FreeSerif 0 0 0 0 VDD
port 5 nsew
flabel metal4 s 2368 4410 2368 4410 0 FreeSerif 0 0 0 0 VDD
port 5 nsew
flabel metal1 s 2623 4788 2623 4788 0 FreeSerif 0 0 0 0 VDD
port 5 nsew
flabel metal4 s 2368 4410 2368 4410 0 FreeSerif 0 0 0 0 VDD
port 5 nsew
flabel metal4 s 2368 4410 2368 4410 0 FreeSerif 0 0 0 0 VDD
port 5 nsew
flabel metal4 s 2368 4410 2368 4410 0 FreeSerif 0 0 0 0 VDD
port 5 nsew
flabel metal1 s 1720 5170 1720 5170 0 FreeSans 480 0 0 0 INN
port 6 nsew
flabel metal1 s 466 5966 466 5966 0 FreeSans 480 0 0 0 OUT
port 7 nsew
<< end >>
