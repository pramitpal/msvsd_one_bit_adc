* SPICE3 file created from /home/pramit/EDA_TOOLS/work/week4/Manual_layout_ring_osc/ring_osc.ext - technology: sky130A

.subckt ring_osc VDD Y GND
X0 a_173_115# Y GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X1 a_173_115# Y VDD w_188_178# sky130_fd_pr__pfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X2 a_312_n12# a_173_115# VDD w_188_178# sky130_fd_pr__pfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X3 a_312_n12# a_173_115# GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X4 Y a_312_n12# VDD w_188_178# sky130_fd_pr__pfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
X5 Y a_312_n12# GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.1218 ps=1.42 w=0.42 l=0.15
C0 a_312_n12# w_188_178# 0.09fF
C1 GND a_173_115# 0.19fF
C2 VDD w_188_178# 0.15fF
C3 GND Y 0.13fF
C4 GND a_312_n12# 0.18fF
C5 a_173_115# Y 0.12fF
C6 a_312_n12# a_173_115# 0.08fF
C7 GND VDD 0.05fF
C8 GND w_188_178# 0.02fF
C9 a_312_n12# Y 0.10fF
C10 VDD a_173_115# 0.18fF
C11 a_173_115# w_188_178# 0.10fF
C12 VDD Y 0.12fF
C13 a_312_n12# VDD 0.17fF
C14 Y w_188_178# 0.10fF
C15 a_312_n12# VSUBS 0.23fF
C16 w_188_178# VSUBS 0.40fF 
C17 a_173_115# VSUBS 0.21fF 
C18 GND VSUBS 0.01fF
C19 Y VSUBS 0.60fF
.ends

.lib /home/pramit/EDA_TOOLS/skywater-pdk/libraries/sky130_fd_pr/latest/models/sky130.lib.spice tt
X1 VDD Y GND ring_osc
V1 VDD GND 1.8

.tran 10p 2n
.save all

.control
  run
  plot y
.endc

